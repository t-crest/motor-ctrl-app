��/  W�� Օ{���.Ebpk�Ǚp�w=����'_Əyka]�Z���`]@� *P�RÏ�Q��P��o�v�Sֈ����և�x|���c-k��\^=m�����R*~�ؤ;����|�f*8�]���=q�XWuX��y7�<E��z��K�B⏱h�v�:�� ���X"7[m�.w�rApX��E��l/�o�3NȽ��oʋ&��B���Oq��Bz��KG8r���F6p[��J����(��2ʺ�g7�_%��'"��S�~{H���%�5�.�e(9�ܤ����đH8�v�bp���j���@��A�9|���!�Ӱ����S��L�r�٥"�G�ۯM�#���c�V�uΓ��׿1|	�0���̵�8`;(UTh����Z���=�ߑ=�����c��իI=uyN�w�!��z�0�Y��0z��9c�`��t�6���5Yߴ���KM� ��x�긾���I�j���Si����!�|�Bjâ<�K��e>F���il;]�զf���/v��Bf�f���9z���Q8Xq3���"�y��c�=���P��㧥��N���:��ү{ʨ��_D �&�:5:XdL,]����'09��#�T��Rm1��,�hg�H��R�e�
S���i�>��|y˸�<�Z	��:Cf�Qm�"�li'p<m�Y��d�f5�I�z�O�:n�=�#	�ZB�5�N���|_�(Zf�ԇ����7H����2I=&�C�)����k�����9�J��[:����-�9�qh�@0,]~���J/g9��\3��/g�K��1h���z����łUj��˚��A�eoeR���J�=� Ֆ��겛7!���2���.SǏw]��D�oHy��$��w6I[(p7�����W��VJ���ҧ8�Qv*O2 >�p�ِ�!����`� d�ג��P�9�dd���5F
����P�b���ffe��>'�萸��]j?p��l��7Lm}������l��Y* �ȀP�T�������tҍ =��K�~�Ϭ��#Al������3q�9CՊ_�M��=M�5ZƮ���=�!~���6���,�(�@�.ԟ<��g3���H��R	�Y��[�E��@�$�5`��������!<c����.{?t�C���$M�G�q�3�܁�蟩�p2�/����8������Z��O28I,���.|D��5���� �s���T8��a��=����8v��7�S��}��F菢�@���S""��Ay���ovO�{��!M��"]�Ύ�od���Cͯb���,���,�M���y�	nȵbC2�l��V'0��*��[���
��vڂ�mj]��Y����W� ��J�!�[�Yb��ZR�3���.X4��9d��K����������Τ�{�������=.��,��� �m��l�P7�ƭ�".�|���R��:��,qKx4���wm��Ɨ��gd��w&}��t5��8�?�qӿ�������u�}b�r���T�~~bQ��?	�E�����p���ȥ��k�T��.{%�B�v����-Ա��?��~��t���ր(�d��h'�Й%�0 ������a�6��t�5�/��Csn��D%ͧ��9��b�ڸ6'FF�k�J�n3.eIĒZs C�בQ�ౙ8�1�E�⚎`40�����ǻ� ��w��2`�4�оOq��L�<�tj��[[N|FBiN jR?l;8(=h#Şӥ�M���ׇ�v���Ɂ��z��Ź�;���ϱ��<�o�`䍵���.}?7�P4g��D2�S,�/�\l�̱52r��%�wq���i�L8�ȟ�g ��lz�,�z(ywtV�/�8):ҩ���KH�P�l~W+�$�L���t���m-�X������KzXE�x�y��[J׊e�~~��qa�bo;���֙ȧP'�pݩ����b��Y�a��,�5)����O7��ɣ�}4�l�_W���ygR��s�Y$��v9�!\�c2$�w6L�/˜���8��%���� rM���w>��%�%�F�"B§��Oi�M�t���Z�X�^ۓ��𱄢e~��f�(�ѩD�X����g����-B�}�)�l�Ѫ�'�ly(Qa��f�#|�NJ�|x"Yq����`g>�A�R!��F�ϲ{9j�n�©+�3sz��#^�G��$?�{�8����\�Jۜ��ϕF��W�_3 Y���&��UcA��S��ȗ%{Fo"֪Hu�����hcȦDS�Sh��j��̭pm��`Y;�,<�{?f�&�2@=�bh���#��#~��\IY�����TT�Ш�S��ՀV�=�W��53/#j75�u�������nj�,OE��1{J�a��7/� �;Ҽ1!(9ا�+�bh{ �0�Z<�Ňe)l��A8���͝���a��M��a(t��cN�ԣ�y��u��o�@����j2 5��Z��{֤�k�V�w�/��ʍ�q�A��e/����(�D	lvPè�����V�
|�$�sZ]�r3��KI^�?t�M�9�`g;�; �6���tc��d��6p#LrYetIߺi��G�zjde�,�����贍���+�>�e��I�'v\=�e!@dW<�+�rq�&ψk,&��B�ȩ���O5q�f`򊨵���Z�^C9����w��>� ��Ny�p��� �¦73]cV�ˋ��¸}R��;c�RƩ���녾vm�ZzڍZҝ$�$gxh;BϹ����~]�v��0�mS*v/��Xd��Ti)w�!���l{�7�Ѝ'��Tv2�뱵t��W��wV@�Z5������aϛםR��|�]$.%�+!�Xl3'�N���"��'���Ȉ<� �^	�}tJ�Cc��]���bB7��_��J���W�T�P�v��8�M���h��b\&��1��Tl�8.��+P�l����-T>X�c���{��E+��V����ъ�Ǒ�>vDt�X��V�}���Y�?6�����N�D��گ*��G�,`C�/X�+�7[��:q�K�yM���� Ul��t��ּfG��\�e�Lɍ��hl"��;���X�x�����i����X���d���]�2���+���*S��302u�(|w��ra����D��WE�J�j���BB:�U�T�ݥ��#ݸt��`'�5�H�v�!KМ���0����֧]�@U6�AK��ɔ��n6�h ��壠�Dv�� '�Kw����Rp�hh"��`ﴜfyX��E�	U�V�	�#�x���S:R�df�˜*"�	g�)��� ����Qs"�pZYv�&�g��(��jIG�j�F���B��.���6��5M���%�R#���6���&�i	B�"�٢=Բ,+^_A��3`m�߸��s�i�ø4Cv'�ʨ��8�-��E������%��K��K����z��q���$��o]�E4�:d�0�Le�3�E)9�R�6>84ԅ� ѫ��J�޲E��,�Blp�L�&]ah�p��e��[E
�����Q֗�"�ԼA��؝IZ�(�{_c��<|���\,��\Q?����(�I������}�Z�[��Pk���m��`8�'�۱���-a�^�u_��7|P	��˨�"�;��R-@��!^�y0���W+����f����m�$�� ?a
�c �2.�YSy����I5����a�����fI�-���'�L��6ƎRF��>�js����9I������<��ٓ��rc��*n�[s��|�5��_����UUPRl��\��n[�]�l��`�zG�Qu,��p���>ÀR�ХgU+��3�,�'���X^rps�,h�x���@���[�7Li��N�!#;�4�eQ�h�E��d�6{�O��Pbv�r���V�B���ؼ���X6��*�P��)�z��8
�ePC�e;�~��	,�wy��`5*X�c|dy�9Z(/�� �9!�q�0�� >����}�Q��5�+	����"n����ek�]=��N��������ͪl�p.��,X�'��<�M��{���^5��0"����z��I�3�b��m��8�^��u�c��0�`�� ��b�1��[�-�nVH
�W�mnZѝ�{��k#)7<7g�q�A��M�}�u�6��4������#x�?1&<E/t`�Iq�=d«��l!V('�ǃ��@��_��Y�1���_�IdW6��&��q�,v����p�[�7���d�����\���/�y#I�e���e�ɒS���~eY*�[3�r x�Z�ѳT����
p�p�R)vM��Ԏ�Ǯd�꺙n6�scԁ�>#�m��F�x�HU��y J.�z������Kп��~2��r�9�4�0N����**�N�-�p�o�-���z��C�FJ��2�hJF7ʬ���
K-��ց�+�~=��߯�Sŗ���"�r���zE2EN ��c�o��6��Mx��0���OG�8DL�NDc7��0� �ɵ���LQ��;�`HR�BձQ�锍ދh��2�v�B���m��R���˳��z����u�Ɛ*N���5#�)yq&-C�������i�wu�[���UZT>����r�4�J���Nwj�������a�z��e��`T*�(
X4�����kE7��.�#��c���VV��u��]��i
D*�V�	|�UW�@���Ŝ���Q���#�}�%G�/�hڢ�D@q��x�=Y�E�>��N�b��@xj�(DS!�/�Z��kpk��:�x*��q��?'b�����������4!��A2C���?�&���[�ֹ�	�y��2Ţ�9ʠ8�b�����*IG|5`W$�X<n��>�a�L���Q�c�i[K�J�)8]��:���sM�e��� "����تuj��#�d��Қhe����O��5������i��4�P�~0�Uo<�%%;��Т��,7��#e���I;H2����h��b�s&NШ��8�(b�F�S�L�����L�h�g�y�[[��	������9����E��!޶�SG�a�,k�86I
�\��_]�t���3>(.|��&���Y�@�_�����^�|�^�R�~����ZB*�u���F�a�z��섌��C��	��k+��5���"x���h�Jl�KM�w�5\�B�!kcA�=�+���4]�Z��k{Aj�c���A�=Հ�~����f5�&_���ě_iO��B�J�[yRnA�`x� 0  ��(�;F�AΩ6�Gb�
髞�aG�C��8T�߬��ܹmS�0�c[|/x���ρB78�� �6�hj�3c?����)�b�*N$��'0�xC��9���-������׷��W9i���`��Q�<�,0�A�D�!�v�D("H��<���F�	���ji��#��]��ӗ�.0�~Y�^�,i��壒�q�07��De����K�3��D��� r%ɔ��'t ^Q	��dB�9	���N�U�XR��cݔ���D�n��V�컕�|�����O�ƨMm�?IY�t�?N�_�{~I���rj_�[�@�-н�5"�����b�Tr^�q)A�7�E�(�t�X8敺aU��n�C�֡�^sH�#"MFv�QW�#��d�br��� |��C�z��v�b;�c�eJz��� ^	�%�x~��ٽ�R3��W��I�X��B�'W�L�:��L׵�K�Q�Զ��&�9%q�1�a"��_���I|Ɍ���6�G��!.
�ƾ5����:N�M"+p4(��Ү�� �0!%�a�q�Ͷ��z�����z�DRY��^�W�w̓bN�hc��B�ӯx�f=�<���0)���T�T�(�^���"�F��O+A$�i���F<L�<�ҙ�>[�6�zy�x+�s�Dt��M�Ĩ4{`Xw+��3;p�T�v���?���|7��E��nJ�fZeM퉜�	�=���NI��:^���86��Ɓy�H�<�..ԘE��֘��y)�q��.�r�$61oO�d˓�dXX$�����s���`���?;M�^r�r:������:��52��'�1���js`!�y��[BT��Z^ߣ�
#F5�z������
�WQk ��u4�!���x�'��&��;&_��V���Lʩ9��S;M�rl��/���+��㰀�F�!	O�i��k�9_��&��]���RU^F��OL��h�E����:�H �&���������ۢ/����C�2�/�2�g!����n��QW�兰u�0���s�\�dƇ��si�%BE�5�-^�����u�t�[N�[C�N`�MF�M�Y�<"a�E��iX��t�_NR.���%d��J����+��tZD�>��X����k۔LA�P��	�@�����8ƍ@�)��:�BpbU�4c�`-��*��d[��}jהc�&WuGu���,e�2t�^�jK��J�i�a�� �_�]��./	��V��9=\����o�M ��gem{�A	ξZ�m�����i!�g��/A��W���<ǌu�kPq�4	�K��|�/�����T�������[��Ʀ�U
ׄ��e7�-��ߢ�<���P�o��e���jX��ู�X�l���I���+��,�:P�[H�y��x���v�`��d�@AӦ%�p��mL���#�%X�BJ9Wb� �EE-�/9�J������e+Cf�i~h0!w����F�H?]^Lb���Żf0j?��l3��t��w����t:���<xO��Ղ�ɫ�(���u�G������Bz��V���ش?n����oa$�Q�j�Fap�K���Ⱦ?F�[}�H�Ϡ�$�t��s��$b��M��r~����<�V��V�)M5��4K��6�(��>e��� be�r�d��x�&wD�����-.i,6�s�_k�6�H2��8Zs'C���IW�s��NW39>6�zm�A�t��ѯa[�)��][2NC��c,ȇM;�<ŋdF=;_�5�n���}j��4i�a^���y�t��g�87�~�!