��/  ��>4=�}n�Ma�"�[�E=q�qO�	�g<Rz����.�V�IU^�G�9wN����-�N�O�א����[�yp�&D�1�Y:�s���z��g*�y���՟�￸����L !�uk0(�Q���ϰ��&�&`�4¹��y�K���(��cɼ�#;�^��<�J���6�����֕��**�4�`74$�xe�#]k�<DT�=�� �M�-ΓS����H+��}0�F�]���݂���������(4�l���5B6�A/�>��0h��>� ֠��Q�5z�I�r�8q�+U��?F83�?c0�<�|����y�am9�R�˩n
JƸ��t����l=�/�J��G�lR.9:�	���֧� ����䈜&
x.��u8��p!G�����U�S�ӥ��}l��J�6�~Z1M��f6�R����(zb����)z~M&K$wnm{�v/�Bl,D���D�q�V��.�	t��$������^��y�W���"1�Y U���o�R���h�0��R�5����r�Ğ���3�]�<8���P�<�ŷ�oB���u�?XWȞsĥ��U�>C������d�����k�)C����e��2"�g�"�
�_;�g{�2��M��
p� ��ܓY�*����ݦ4.�ӹ���F�2�s�V:�1@�6�F�o( �"�^d�&�P�<A}���/a�A$̔��xuò|Cz����b�l�y�Q�j`�c4�L�<�8��AH�/l)Ҥ���ΩZ�堤�EZ(*�@�m�{<�x����x �K-�Dkc�"O����� ��Ok�|��o�d�R������y�jP��Ey�<D՜*N�֬�)�1��X�1�A� {�s:	&�}�=��]�{�ŉ=�ѐ��);dK �z-n���(��	X E{¸���J����S�IE����$/1��v��f���U�IK�Ua��`�M���v�Aw�*�k�8�7��"�?�_��OչGP�Cc��g�DW��H䨬^Rh���j�P���Tm���F��򨂘��ef�g�&T�Ĝ���~�\�xʷ�`Mf��*��9δ�V3Xg�2�76E��W1r��^)\3���b����*4�O�K���`8��ԥ�� ��f|[t���8���p��؉�i�x�Oz�\�R�Z��Ѥ�rHH�EOO���@�߀>�GA�um��D�A��,eM~��oB\���ݡ�e��je`X��o��������0+�U ��$%�ݮmQ�8��~�)��h�{T-�l	��rHʼE��t��q��d\� Q�D�+tU���h��~5���E�2R�&H�=��O���A�oK�[�0������2?�|���_�p�E������Yv|{��*d2�L�R�a���ap�O���%٠�4r����ԤQ��ʐ}yʹe�Hr-�u�N!ѕ�<zDN �ѺB��)�E#0���w$1'�'t������'�8�֭Z��쬰O�A�V��$rG����*{��
%\�|rf�N~1V��A�\jJE����3Ö��L �"
z���r���h�e���ǂ5 �bу���Do������Jx��ʄ�WO�0	�k��f�㥼#��p��n�	�� "7I�5�@�*�����]4ا�Jd���z,���"��
��A�H�l�.�$�H�5�?i֧�NVw��d�ag9����k@��x5J>q3�nC>P]��F���a�R
�߳M�Ƿ���E������3�mf�Ƨ@��� ���9�ϧ��E���.P�a��׸��DIʪ�QMҒ����G3�Z ���O3d>�/I7�u��%=Y� \��W��4�
N��̇���z���:��*�+����p]������r���$���� &��GzL~W���VL#B49���"�Bg���g�A�L��M_�7̍,Z*܉�4+��ضZ0��OXH'}��Rb���XL�Y�j����;����n��k�B����lg��aZ��_z"������䐜�"�,h�DS�x^�}1N�����U��`l����]�,35ױt=�;RX���$ߩ�}<�R[�#�:VU`�=K�=����Zx��$S=�6�q�dLt�.�6+�@U��ҟ3C�{�z(]���0���Rh����U=�c��=݇q��f���m�Q
��z��ꈱ�-��}ڒ�T%g�a��ۯ	�@@9��d�oJ�R��EW��o��;Ox����Gg�2
�`j���2�e����Q2��랭�)�_���BO��č���1��5!�
|p��00{!������E�����Ԧ�fHKm=ZF
WJc��tr����b��l��?[=�:�e���z@�H�k����Vv�!�6���:�%�Թ}+$H���@2i����d�pWt�k�yHL�yioZ7�0�(���e`=j�XNuQd�����>�:z<s*F�y�2F�~����2�S�O�Ăջ#���~�#\iӓp'�e���{#u����&JTS�`f?R�eO*��QK%�~p/��?cXQ�(�p��"^�W"�&!�=p==�@���]��_T��^J��b]Y���r�ȋ�.9�v�z#*(�#��<���e�� ���|[X�Ǜ�{6��JP�cn9cI$���Y�w&��ݼd�8ӹ��iB�cOR�'���\Q4l�ߖ1����M��v�aό�)m�%�d� �ޯ�O��?,|��^��d�K��u_�F�ΚW'ȣ�P�{�j�)Ur��x��3J�V��,�g{���LO�h���.�^��z2%��A^�	�/C_�X.�%�-j�_��������h �(_�!Z#Aͅ�Ȑӄd>���ݤ $�\�nk��πk��3/�D�3��8��:�f����h��R�.Z���`�&�P�����.փ�c=�L�d,)����D�d{fю܋��>'Cv�Ϸ�e;�K� ɏ�]�	?�W�яV9��~����l�3%��o��fHqĕ5zJ�/�ZyB���,���5��'y��)�fӵ���h5�V�)I�0w(E� ��"(�ٲ�d^AN|���q~\ud:_��dp8��r�/v�G���К��2a?$W��U-"�.���_zBDI/�:!0�շ���� �=��z���epg�\�W� �:ӓ�5^�I�Z0T���V�uL�����1N,�,k@�5�Տ�D�WiY����ʡ���3y�b��CrD� �$6�[���.��
A��Z�0	θJ�z��!��q��z���S�a�CfJ�E4q�H8y���ٜNY6ot����ɬ�I��8S�+�k8w���P����c�'��R/�mW�/ܨ���pe\W[�E	������F�b|�jn�!
���Q�:������ؗ8qT���m��{�&�@���1*��&���נ+m��8\M��5:���OԻz�<�K�h=�P��9��.�S��p�}����I���%}�Z�%tM���ϣ�җ�fz:�PV�Av�4�P�2\&w�Gت@0Y�m6!�6��� `U�l
���%cm�*cx�(��؇���iM_E����"`Ālq����\u z4��A��1�_�pኳj�%\߯�h`i� ��E}���Hk�E�C����x�+ldES������BP�8���)�ǼЍ�@A5�P�^�j�������1[������!e6���/|�ox����|xl?��>��ڪ!#�����Mٌ]ى��������U;��pHK�o��e\��O��$��RK�[*�}��@r����$���_��\(c�ƭ�s��by#޸@5%�U}��4 �	��P�W\�x5b�i�����oLlk�J��Ly./��P�'�y�^Kq�z-������W�W5���9.�cQ3�
fײT�o�B~ֵ%���'�����yF�މf��!ߗ.�_~a@��8k:���S�T���	�����Z
c�n��v{����>�IXc�H�FKb�*���E��kp�B����{L9B���f�g�����}����ˠ����j��l��2��BA���O�C��%CXC&����]Ɉ\D���C/�u��=�2�Cg��e^����o̒���f����A�Z��n0��'��;�7�J��ا�X�R��M4h��Ϳ٤����*Ř!�:SH�.�|�Q���X�(TK���X@a�;�IHBӫ?�"�a�G�g�4�^�`�3��>6:��t�7��.�,�]^Bzf�����É���Y4�j��>����n3F�Z��_K�D��:�Uq����	��}n\�"˵�ֳ`�ƫe|�u+��(��ʎ��-����
�%��+W컑��yj
.f�D���!�$d���|\6,�,������҇"�gLJ�%�ͪ3>�B(yü���W{�����F�e��<�}�e���%���������]}]h\�ڊ��3��O]�q��R��^�)c?)�_~,tx2�����=j(߿K�	�4H�;p��9�a|O�CH������C*��X4�R�mzW��¡H����$y|����].��Os��U�5P%�dd��0�2#�w({Og�����] ���ef�Z��N.D9�������}_[.�S�2o��m!=mū
<j�zTG�O��x�~�u�.>Y�Hp����Y�� ���Mգ��Tm�� W�CG���C+���ԭ_�>�1����P��!��Y�r�	������f5��dg1��\͙�0�U���H&
q4;�G�r���Bո�)��0��00/Ufg�_��(Y����R��=�X�J¹k:|n Sa"�ڼW}�)�Ѽ���-��d����lh��ᴱ����SN��"��2�L}�j�4p�1�q�P���|��p�;�H׼z01���f'$?lj*	Y�|z�B`?߻��}6�_b�wH��C� X�Wƅ�+���h�y���Gg��l�F�Vd����W��b~{�O[R����w(�@�C:娟@r��<��ʌ#5 q)r��V���m�3�@�6�?SJR�VA�"�"�U�0�A��^�qEHE=�ޏ>���f��j�oOR�E@��We�IR�_����9�|%�u��j�x,k��(�- $<Z-���fֲm/�%��V�4'�e�Y��PEo����r�L��?�GQ�A�c��k#�I�t�@�H �~��K , �uM:7��5ȷ+8-����]���Ug$������ItzfdX����� ��N�[��MK���������/ A���|��.l�F�-�B�:`�(��>M��@Z�"�8�i�rA�z���XI\�2'��K��%���0 D-�~S���@{��Q�vX)��1��"a��&��GZv�%:�Q�����aV��!Î��\�����yYD�����:fH��	����u�Fs�&i�O�ŖNgl��jFa��k:��S����(�����r�����|���e�Dq'����	P�M���Y
��e��� V@��wA�w���k���̦-�6�t-.w��mp�S�/�]�ȕWh*o��֎����YC�+	0�>�>�{{�	ư?�p�,>F��ߴQ�O�^P(R'9�����}����JL�mb	�J�����v!�W�c-H�'�_sʾq�̣��'S��=��5���_�'���m��|�g\N�Z@2�Ru1�5ć�}��[;��,�����ٌ�i���,«]M'��Y��V���>��ӮWv�N�lY��/��a�^\��.�M���vT�[l�h1B'���U�C��X�:,��4'x[G ���q������-9�K&X=��M�\�d��ѓ>�}5��D��+.2�f��}��P>��������6t��}�2��u�"e�%A����@��1���6K�jH\�de�؏Z6'2�=�$?�O��,�u[#��er���R&-�bn�;�e��>Ӛl.D���mO��RUJR��#}qf�	���+a���Z���}��r�a��uL�m�&����JjJ�U#���ҹDK���?t/���\�o�X�G��K�Jl�����w�k�sC�ݶ;\<y F�{�ubA܈}G类o��,��|�%�|,���dTD���[@}��J���͸�=d2��y<+ �~p�'�Ҏ�\��%s��o	d�$����Z��Y��6*�T�Wj��y���:嗩ݜ0OJROu� �֢�/}��n:�k��!s@��ٮ����zJ�ePT�F���o��}�\fk#jx+�X�������O�9a-l�q`^'���ً��0�����f��P����]٠����]��#Y�c�q����}G�1�`��/{h�B�[|�$�ǒ���|������+�	��t���8�l`�6.?N/C��u�e��r}�!��:}����i�9��.�ĮE�����?�s�7��qz�Ej�c-x������?⭦�Q`�oؑ�H�DY�sd�0yZ��n���^>F`o����0��8�;���xzWn��L�W|Re^�F����=&4�V?�!���(7�������^�ϫ���>��:�?�v���T�Ok��)J��Z�(@�E�H��
�W�<˕"+YU5��M8����b������r������H;���Iv����K�Y��.�!�q���� �W�R�?h���b����Kk���%%gs������o��QY䍕�� ����=*�j�җ��_u�|�D�Q]6'EÏm����y�B�6��>���X�Y��b���A����xl�n��w�����N,Xt�:>SZ���� W����3�=�tJ*��Q����8=��e�1��޹��>�3>��6H�f���LSi/�w����ض������{�?D�t�g�G��χ�=���J��>�J���m��Q9bs��37���_�H�*�^�H�d��E��<	}8=�p|�n0z�y�m�&�����NGYG���8�
�{��3�Ӳ��S8GU�\D�i�;~DHr>A�B�!R�5R���<Q�[:���R�;�~3�
UH�6�~���:�� ]_� ������������{��u�]�Ӂrq������db�� ����ntu�-���H+��C�����a3n��P9u>[�z-a���oF�vm�$TI�q�YY�3rCHĊ��+���H`� "')>_��_��T-hD�ѷ)چTsB�LO���i�dC���@�I�UHg�O���~)�l"q)=wK�m�D�ѡ;t�KH�����hR�2�y�x��d�~�ndզ��{��7:����xkʈ;��+"Q^f}���.Yu����R��� ��1�����,���m���랶�b��®��'�^�C�	0�ÿq���� ���i4�3��u���I��*!�||�ݾ�#3���/�iIJ�#P�d�_F]�mkCp���XJ�����JA�%��,)�mb�����G]�)�F�w�[~��o�0#{��z��:�͏��4}XO�{�!G^~�}4�����R3/*� �Q�u���!�L]<�q??c��� T�T�I�z��) UH����ʞ@d\������-C*�u�(���@�-��c�`��N���G��P�ya+aG�f����I�C�ܸ����3oH�vIC��x.+"�ͷ����}��s�$v�6Ƹ�}��,7TiI�
%�^����He��OT�
��@��+�!ɀ�^i�$,?���=����Ħ�'����6��Ռ�i���I�W���:�Tg�#E4ۧ7�	��]\�7��&��D��E�1W ��x~Ʈ���I�-�o盹�0�UӀ�%��o�xV����'��F&ǈ�����V�
�	�F��BC���m�)e4H��@?�X����B/ sEc�Y�^���� ��t�y�ŘU�� 4V�&��"��GB�̀ �K��d�� B��~'��s]������h��������*g` e�O&U|\�����t>�\��1�2���+f�g��-���K�B]@)ϵO��+���������'UR`�m��b,m)H_�b+z[8����l#���u�>54���9�vx*~���8s-.��$9٬ø�̏|�A����Fϥ���-b���MԼ�{���� �Dr�l��k��2W�/�)���x�����ץK��ѝ�+�~���9�Ms��UJ������*D�S��^�@ 3ai��
OJ�[��K��\�z干NSIz��\.O���(N5^��W�,���{	���������W��,�߿�.�?�xޒ9T��#�,$�R\���}�G��|��=�����+�S��n�ZIHH�*~��:�:8$�"6��T��='�ᔖ�#{Ϲ��=J7��z8j���A>0��ME��e�����v���{��|�ޟ���e���d��ޛ6��$&�҅�c�0L�����WC�� TyU����peCv�܅�7ʺ�D��!��'���H��b&Lgb��;D�������b4<�O��O�"W��ʄ*�[�����Gy�&<4��{��O��ӜCl��
e���u�D4-����na��-�՚v�0/�w+�¯gl�����ʾ�8X"�0���J;��f0Ih�=��VN��P��}����n�]���rTL��7��]�����{�S7Xu�#�Z�iȑP���>AL���I��HB�)��y`��kQ)���Cy8*�s)�4� ��	���W��q��t7A��˖��=YǷs�ͥ]�^�p}eyy@u��K��O��A�S��h&8����@��?s'.8�g1|q�v�f���c8����CB��70xu�9 ��H�iUu>K&&dI{$A�u*Z��A��nar��<\T�|(g~Q`�b������p��{D��|�A�ҀV�*O�D���|K�0Đ�����~)GL��b'�%��u�LHv��Y�U3�k�q��_���i�ksk��%Z�v%%
X9���n��qZ	��
�+4P�^)�8��KS�k��������A=�=B��<�o��),�m��H�E�!�4�G̕Hԭ^�����i(QG��7K�BaA1���p�����qn�,Kg��fA�i�s���wr�R1�x�>F7�1���>S馜C�5�t_A�n�9�����L9=#��<�O7M���ǡ|��o���"T�&�X�|���>�x��y�(1�Y8��)���j����h�w�t�O���ܻf���s�tU��QH��Y��'w�⑹2�ʏ�ud�^�d�r]k�'F�KYc*!�>��r+��^�*��lMG9a_M�;���NI���P7��C����6z�4�+]C�Z,�kT��7�F����ޭi4� S�,"�K	*1k��W*j��5[QNKo"��(�w4_��|m�k����m���>����/��2� ���2á ���<��R����l �SW(fB��?jH��"'O@5���(�w���� Ғ�\�֡�ڎ����!�������үgX/�3�8���-�Bf�8�%S�O7��Ͻ����5��<�k���j"{���f
H�S)���Y'|>��=5��^�'�8>P&j�h�������R0Ѣ`_2�0?�6�� 1�hR�=ظ�K����d!e�3��m�ϛ��4d��V�p*�6��i��]�
&v� _j�-��#Y^�Ux��B�9�5+�n��^�ɋ��J�$�v������-Ũ|�Z&;5��T��\,�cB[��1�_�H�wd�c�%�f]��o.���Ǎ�	�h�N��N��KEDJ\@i�戈p*~���v��)�Xi���Cn��T�}'WU�7��47ۍ�t���F�&�]tα)�pG��n˧��Kv���TKT!^).*��Je��O\ݯ}e��$�XH���d��{���J��R7���5!�2q�gbν��=�k`��Ϯ�ǅr@T�_ɦ��:N�?�c(�k�����9���ArC��.� ��T<VR3I�i���j��A��$c^�Ӄ)�6�0���b�Lw'*Y ��3+�Sۮ�����?i�+9e�>���/����K��ZC�Z%�� e�W��yd/�w���~�Fu�6��AT���(�D�X?���J�O��8�z6����]]�K�e��wܳm�u�*ݡ��A�)nq/aP��M�F�a��p�JK[t$C�f1X	�����+ #q��r�n1Y���+�!�-[V�&lZY�DN qe��t����h����ieZJ<����V#K��w��A�9KY�D��E*[ ��s��*0D���O4���Qfe �;�jc!�+C誷���s���QA��;]"�����2S�ԗ���A�G�5�1�(���V��m�	�,�#2S�,Po_�! ���z��%��&�?G��cj,k�����4j9�ja"�������B��6-�75��u�ˋ���v|yf¨N�J.��"�y�N��R�Bj���b�XZ)�C�K�$�+�;��4N>��z��
�z�V�e�X^K�%e�p�����}e$�!�vXfq����fd%B����w��Z��ϝ�݊�{pZ��҆�ꚢ-k����j�蛹M�� �9G�$u�P�v�B�e�x�H&��:�����l�����,�����R��#O$1v��� �2���^�5��)ѵO�
�Mѵ_���(�N����&�XY6�;>J�<��M���u�g�󘋹��&�rdb�>nNg��<�1��ƺ<j��ݖ4��53�÷����A|��f�����U��F:ŜE�&�y�.�&���bݝ$`ځ13�D9�E�B"4l�5�ԙ�T�&��P�3�E����_d�
:�  �cǣ�&��⁉U�ֱF4�j�Qf�s���%O�r������'	B�m�����9Ϸ�jj�ǧ��;�4�}���g�u��*C|jFd���"z���k�@P`P��s�k�X2G�b�� .<|�+���*.~(�Ɉ�>O���SO��	R�M�;H�L��J:��gdZ�883y>�U�u��)$$�fΨj�Ad���7$s���(k�w�ֳ.\L�V&Zb df�]W��_$-^ϸlAv���KZ�dx֡F!،Ŀ����;��m@b} Ѯw����s��Y�ǥ�x
�*uH¶����oE˽Q��ƯekY���"=�O-Kz6w�$.E܉�%�7���� rfw�Z�}K�<Z�`MaT:�]�7���a��R�CQR��&NMlH���Id{p���/y%v�Y�ٝ��1"����x���6�F8ؿ"<�\�Di��03��4p�?>ޯ^�栽�9�$6k-�y�a�&=źB=!�^%xx�p�Q15���Tn�雚��%E,s 	?�-1��U���T#L�x�"�������+%k,���+��m�VΎ!;�k��~��8;_b
�AH�ÿ�����ҥ�W�}�
=���V2��lTC�����Ƚ���|� v�_L�����j����=�OO�95V���3�,mvL�E�E���H�(�����u��܉Ơ睰�&d�y��6��P�����ɓ%�OZ�>?�:J���i����/�����Ĩ���8�y�@�|F�GW���ƞ5��#�X3�~���N��5�4-���B,���yT�Y8fa$w���8�dx��䦥lW��1��)�զHxN�HC)���h��p��:øÏ�J���\{E�50�K!}�F��:���p�����`´��Ă�.RİP��)�U�{bkV�"8�R����fW?1Q
��p-�>i=���Q�mJ6Y��!��^R�Ft�^�+�b�a~gBK-b�+�B�W�Y3I;Qpa�V2y�3X�tΗ$o�M����apI��SpI�}%h/���ڥ�[��S�/YV��"�L����D�g����r}�����-`�0��$�L]�WK��� ,�-��v�_j���C�u'�B�ڝҿV��BG.4{��X��7�?��{t¶����9��]wQi�pL�˞^NG|��02R�~�U���1\�N�������&^n�d�~kJ�~ح��hP�'�ڻX��@,ÁU��*%�͞�_���͘	��U�xj�?���Em�
������-���m�A���^<k"��<�+�� v�:�2)�G��-]�.%߷���	#G��;bp�0��h��
@#���۸�w�<��!�:���Ga�Am����Ui�{\�#����L��VGL�@�>>;�jW(#�E��U�u3�U�t^��薶;n�R�����y�iJ8�迳0�pO |�|��"ܟ ����;��R
�u��Ubo�3���
���w`48
����T��\�W���L�ST���^�[�P�Nn�ZEQ�%M⧱Dӿc�ɣs
��<�
����4H	:O��l�ƾ8���@��/\�mlJ�Xk֪Nɨw2�t�)70��gq