��/  ���Kg�DoҀ�X��ry�4�#b�z�q}��b[���b�Ή��@�ϱ�a�ٱ�l �In7:-�M^����/�H���O��#8�;��P���8�)����Bh�ݘ�B�����w��\�ɻ�V9*2�w�����*F��1�a�{/��g!��wU^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK ����E�U,R�v����RGa�z}�Zے-�h2Fj��5�!��k��vM�8y����Β�S�����W:��NNo�?�ݸ�{�qǎ�DR/�iM�"R$�w�-V �U�4���r�O�S�M���S�07���>E�u�����s�2>
���)������꭪�P�#�UoOv��N()��~��o5�BtO�Q���@^�Ao��)�wA��u̎�n�������X}� >�H�]Q�T�^�t=:e�4��hH{�2��J���Ӈ��,ۘ3��Ib��p/�ï3�8<<�ΙF]���nDS�����,۔A@��J�Κ~D�d<�Ϳȟ	�$�.�d��Z������v��*^Cs�Z+&�T��\�Q��=�ג����{���lD'��|2�Bm�S\���i��LM���Po��q�v���CVc�ЬF/7��aT�}��λ;�ٚ�c��V�wQ���A(�B�����H7~��7���o��xH�k��:�A�81�!�Nc �Eq�����|)�VG�L���X,� 	�����b*ᢡC����:�_S�j���8�=��3�~a��:7\MN�Д�:��Q3�/\kez�A+'k�c~�
AN]�S��;��99}ƁC� D?6*�� ��z�toW9b��u���-�j�|a����B�k��Kr`"��G�c��u��{�7��Z���ɞ#�-GDQ��yuS��[#,MH�,�}��"* :��-Gv��T�6����{$B��Jq��g1��eˌ�T�Y��t-�4�*����,�tI�����<�sn5�����rq}�^���D]�ӿ!p��'���p���$0�c��}YN�8n8֚�1��N����-�f��7+%bu�w��t1��Fٿ�ne�-�4�L��g���d<��<���#V� yfyE