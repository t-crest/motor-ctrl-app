��/  Z�OUEZ4�uZ���cTD��[���6	w;��F(0l��$��`6�-�2�+��7���? ^���j#m;%z�4�T}l��@=���d�Q���۝�m�9�(�����7!@{N�G����߅�=�%%��+~=)��uZN�įdb([�l�SSM"��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<v�d+vw.����M�ߖ�{���)ٰҴ���V����-�x�M���`	�/���B�O�Yh���B��^��D�S��>)f��4vz�R��6��)���);�ߔ_��*���t.�{P۳*��m��ߦ�ԇ�fL���6����*c<o�1g�����]$T5�G��v����j�$�TM;�b5�_WF8k\7�r�d¸���W�;��O�Gp&�4���dQ��,�^�a?�˝A�����o�a|ł�8!�"%�!(9$�O�"�גdf����g�Z �jI��w8�<F}�9��Q �k����ҥ�_̏���[S�Ȱ_x���q��JԮI���\}z<#_�!����t��L��@��NYY�o���_����D�d��F_��ӂɔ����s��/9I�_Q�Xt'���Dٻ�i4ч�yu������%%���?C�wrI�S,�&m�}|�~_)z�&v��о1+n�C�!NY�����������P�r�@ w93�i;��"e��g�}Zl�(�*�d��l2y:�B'-�<���}՝n2@[%�`Z}(�kf�����8�S[H_t�b�29�"%�IS,���5W�r�P� ,,�l�C���7��ݻ�?{U�	�mUG{ɯ]�]<d�}��:��i,Mf���+.4��j�v���� �����s�[�K����`8����&'}�,��K�����Ի:u��b>T�밆R����U�U�b4J�X�Ȱ�O�~�b^��lh|�_^p1#�����Z翈�6fC�.�f\j�	3�����Sfq���p;��6���M�[���U
i������Lvk�aʃH���*X�^�+[�"��m&T�a��~�"�E;4brl�݇<�i��.���\݇P�C?�G'�d��9U�_�9�jw�����y��A���Hx~�Ad<���|/d�%g!3.�Eݧlc������=��.[��s¯e�D\���J��$�����a��0��Q������':~|�+��­P�u��!Y_]��6�=�� 0������:5mLALܚ��Y>�����,U�I_�=�Mh�M?�{�t��6��H�ܩ�[M��Q��6Ӱ�}��P\P6x�����H���aC��2Z%����{gxp`�a�̡>����x�λ�:�P�l���$���7�:��	�X3hz��M㮌�X9>�/̂L=D���'S�`^��H��h�v���Nv�M\�-�Lî�-���j����&�9�`��Μ� �@�`��T@��3�cM{KC��{�Y6�M��vt�T[*Oj�JO���Ǌ��4*���!�d���..������{�3�h����n�f}T	EgCQ�KIUl��pi��!�h~�Q�Hc����Z�t�ZE붻=`��F��7�a�.	O�������;��p%ye�kqmD½�[�Ȯ��L�xS:�Ú���[�0�l���u�=��>�g�J�c��^iz���S5Pl�1<�H���0c��������0R5-\w���i��� V�;��cʵ=߮ݐd��.[T|�x���3|����&�o8j����I�ms�o|�w�����FP53��I��J��l~Jݠ]&�j�P���≮)�I\U��/�s\�a�Y͛��b���1�|�X�^e����"�Q��nn&�$�m����!���i���B���ڌF:���`<DK�aH�k�kNǪ�\o`ŏ�it��#*����鮜�-jQ�
�#��+*5�����|�������ysϡ�v���C�����s��00@��l	^Ë:>��;�����uk(icux����Q-�?�g�L�n^���]���!����v����+/�}�H?�}0�Uíoo/���%��윜��É�W�xg���J���,S[.`��^.Pih��?~�(E�EUmD*�+E?�˝ȷ��;+��=�F�j@��#;o'!������o��}��bE����˔��o1ue0X��G�X�m��$Z����+�{����ɜe�FoA�i��E�ax�����д0=�4�\�� �~wOT)l�C��1�/�}Gpma}g���K��y�AMW�\�-�k�=�U�^�c:�c��;�A���w�����#�0�P����L�In�"�^D�3q�-p=�:���U��ҭ��0ͱ����'�2�2A;m��脩�45���<���"=�#G��jɅ��!�&�<��'��Ty������y��Vs���<<��8&dY�� ��BSk�����>'/��:�>yrEW�!R���zr������{-�v�L��e�gnY6�-��P�z,K]/����[|����,4���lyʌ*ԫ�> ��A����T�n0����*Z�ঞ�����q{jikR@�	��X�0� t-��o��tTs�W!�ׯ��8�a��B�)�+S�+>���c3�!|�k��
^f���]@��t���!������W�n��u�ҋՆW�����}q���x�u�����oƟ�>�%DW#��������%���7|*�]�!��B*N�Z�Փ���:*�_����zN�F��J�Z	U?Y����8f�^��" ������OeL}�6炛��*ܜDh�1�X�h��@����b�a%<hV)�ny)W;�mB�oI=�c��3ɩ���v����3S�K[���>���|t�TV�$�ς��%�C�g&UY�:�3Y�X�izFn���P�y�N��7�9�a��/n��s�ع7�-�Ż��S�(�S�*����G<$OVK�)Y]�`vg��z}���K]�+5��]M���/����㊖�<�}� {LϮ$|J4�l=�U>v��[/��X�XZ9�k�}U2�&�p�,��)�s��*��R��"�}��=b���6������<=���yh�q1�,$���`Q�q����V]����M�`L��!w��9ኲ�K��
��M�U������Q]���q4D��v뷂���l��(��l|����=x-�u�:��^g�lXJV� �ّ�pm���Nt��g�8(���;0M"��"��+3�֋ک0;����-_7Tm*�L!JeV��xH]����>
23E�/��"���8������%b��LN���ƽ�����-�s4�{;�������D�^P�5�MC,����s^�:j��ݨ<!C諈��Qp��p�Ge��ʼ�~�/ޑ�M)I>�U�q� #y��v,1M�%��z�"}&�ay�gOo�&a �;g�,�f�9A�g2M�Ւb� �	ݔ����j�VA�G�ʛW{}L�Gݸ�5m}�pzj��h���ctz�c����,hN٪#���Έ��������!:k�mj��!HY۬`nh������	�-��)\vĚM�c��\5I�ۗiF�5ڇf�ַ��u���կ�ϼ_E�]�$z��r�˅5�-�:C��i+�aK�Ӻ�8�C$�������WSw�6��@~�����n�Q�t���$vw=MQ��nwf����[/'X���\EΒ5װ�����o�ŝ��0� ��]i�U�/B�ׂa�֐�aa7~<�W����K�X*�i�	k�j�Y����a���k�?rj���^mz�Д�L��� �:���ij!��5�Jҫ�`�ێ �������2����N�1�P�2V�,���i�����OH�~o'Wn*ϳ)�,RQ�"�����!v��П�͗���6���`�qC�(�]A�y���^N�M����'x��3m67D�cZAh���I~�0�gIH�OH�-P�H�c�=�{�Q�8��	�O���d�j/���uj�+���Y��*O����ɗT��ƻ┆K�5�L�}!чE�h��10N�H�Q3�~r��B�n�W��NG�o��nF�U����HnK�J.2Ѻ2ʑI{X>f����X�΄����D�5<!A����LK/�/�~b�V<�HM�?�?�}����R �ͭW�����,�3)E��h���1�>��I�@'�e��=�O?	ѧܣh���_�����@�/mœ'2n��B�j�'�������5�~19hSԊ&N�����2�bCr�W2�Y�O����&�ܹ\V�����o8��K��S�ܷ�!Pu!9`TTd׷8�^c*�+���s����?h�2����.�A'���Ҁ�X��
|�.�� �NV���ѣ$+�4�ܢ\�[b�F7rA��ֺR~�iW�6�c�����Z�hµ�{��m{卶��
e������"`X]��A4J��'�������"}j9��NbE �����(�8unH�8@� "��
�H�p�¤���7�$��Ԇ�d�cZ~n&?U�_pY�v���%�)�sd��"9\���ŧ��~=�;���*����b���"D��a�q�R`�B;Í5X@M*ʖ��
�K�/�Q��VE�F����_�VD�~��)�:�g�5&3��Y��[;��P�鴵��h1���<�4�[/��P�0�/b�ͥL�S&���ʏi2�:q�%W� �p��ݚ�V�Z�dbx/8̜���X=�b�����,���d�[.��O}r�U���Pg��ϫ��mTE�'v���p��N�tj�5MB�f.��͐��|�%͎�I�X�h̛]��^X�$"�]����n�ߚ��܀o��A���R��)o
��D�V-#�u�@+L���ĤNU٪�}�n���T]7��Q�����@�Tد9,�Ҧ"�i�;� �1^�
7�)?����<�N���n�M#`�4�E�����s��g���DZ�iX�3þ?')�)w��,$Gi�^�Lj �Ǆ�y����m�}lp�T�H}��f{�q�=�mT�s0!���_��+Q�h����x�(�ǖ�!����ij���P%h'�"�t���u����T|O�K㧮��*ҏ��r߱][iR�����q5yS~��U.S�J�vrK�7�,����q�a��UU��!���֋�v��VSdDvL��q>6�@�%(�s> �U�*cm��
����K\Κ�ί���AzX���K�\W��I��W���������e����'rz�>Q	���1Ќ�.�.�U������÷�{��P@�s���:C_��o��nS"˫��������bW��� mF�Pw�!�R�:���<pS�1s}>=�
�/�����Et(�L��8:%d�VI1�������n����/@'�,����ᅱ�w��z�.�A����!\ڱN�м�%Uh�*�6J�	5p}�yG��%���Z�f��*�֪?���i����+�/5Zcj��/KH*I8�J3v��q�=*_I�i�_�V�.J��e�����xM��L};���|�F���F���lC�jF��gN����C��%e=d���V+�#�>2e�av;����Kb�k��t}e�݉�l��S\�-�$��#��������`�Z�p�Xh���H��B.f��bR��o��Xb���ޘ߿�0�e�:2?�E	>�j;l w�K�+�|��-���9�a�jrAŝ�^0�k�n�V&���2ڍ�h���J��$](�s\~�oY	�rr	����S����
R��Eb��eX�]����<Ml�{��ǽ��fL�{����5�����7�X��9=��a2��k.,�����&��!��EuΔ�� r��?^ۍ�C�9�϶LQ�,���f*�{xݑ�ظVS���F�H�oS���Sp��X���.����d�u�
e����"��}�>��z�Ϋ�"ć�:�x5��n1��f��d�� ���y� ���6����n��?������N7��ѺP N�����I��R�����V����rj�ʂ�x<���A�LXC4	D,�3�����'V����,?����d.�w���F�Ȣ�*#�A��{��ꟳ{g��%��*l)�K�kWa>7��Ɣ��t"�6�(�5�w�z�:
���J�ߩvE�����(�����������L4U� �%G��lk�J~V�[L���V�ܛ.d�`a{�Sw�H�p�;no��V�Υ���x����C���?��d�:���DЗ�����ɪ.dG�`�k
��F�h&ћ9�9v��1�i�ix0�֩���M�v��L�|%��IcL9BM;���Ѧ�;�o������n��y���1��iY�5�Lj�������u��?��V�<�S}Y��D�f�'=F!�Sn#�qE��P���!Ń�1:�(/���F������x^��-rU6�Fo�� A�Q�]R��B�4��p/8ߕP��'	X�ϖ��B�]o��\K\�i}�},E�����Z�3^�2;{U�+%�ULj�I�x��%��$}�� !�B�D�\.�T���~�HG��99E*�(	��pj�~L�x���>F7��ף)��;�*�ğ���\�Ut�8}!!`t����0%�/e�5%D�N}��Z���抍�Qºas�u�p��r\@�T(��|<)6��\.�>_Î"��΄���S�Oȁ��>���Y�|�`�j�[[*]��6�cT6H���#N�>=L^�u�d��/�S���|BĿOe�C`��B;�ZJ��Q�������"YXo��0�c�!�3�_T��������]B�r
�Ș��%lJ�~�ܡ�r�mc����GI���&����0zƓķꮵ�o\�Z1y���w&�g1j��<�t��æ�6Q�$�_x�r�]���w蠡�,CA�O���za�Ӊy��3�U	Z��d�]x�b�$nܫ�l�A$أ�j$�>{;�J
����CH	,>cX��f|f1�k@�'���Ƽ]>�T�j}��7�����!sl��=�{��L-�d�ʗiJ���R�<r�|1���Ptq�^xw֘�_m�`+ֺҎ�����'O��T�Nߒ��X�F�:�q��Xv�#�%p7x�늿K�%�v�"2<�ư�\˓��R#������g��a�dNP�%�7�0KŇp��5{x��v��N�r�����g�8�+�������f[��nl'y��{�\�@���s�����ӂ=�P(�x�Q ��S����]�����A��O����K�z@���B �x4x�VC�Y�	-���wT񚟪�\ B�x�������z���4�z�o���G�T7�i�������������'C0��]!@c�{T�J'gœr�4���M�F���_'�ȁ|�~�#�=��6��L��|/�\�WU*%�c�C���}sr�1n_ �Lew	�Y�{բ!()U����)2X�^����bj�J����oPU(`��VFV���gͰt�+�8��w֏�	!����������ʹ��Dg6ԗ������*}���V� ��S�1�����Mf���+�� ܁���1����=�vE]\���-�v��N�s����%�'�`t�\�H#Ӈ��w��S-j!KX�K�j;=���bڪ��xO$S���ubvuo�ae����!����&��^�0Q�#�)����*7.*��g.6���{X��2���P�e��f��u��.XVl���� ���?7A3����`6ϸ��s�D(M��|��M��W!������$6i4rv��J��c4\�g���F������?�"�֑v�����5G���	����-L����X3�*kD%;�3DA�]�h�Q�-�@�HB}^�4R9\������WF0[acL��Z�" S��z"zk���;D	*�wiJ�l�Ҝ( J�t磣�}��t���������u��mh}��nR�q�Q��P�	��njц����ژ̰�g5�8�B��}�1G#��Ձ�.��P��P�ǡ(8��֡Q����@yD��>O���{�z��yA���<, I*��������0�� Pzb�R�C閱���&�������;��K���q*i��k鼊P.1�쫑U����	�_넬�jpN6��I�Dm9��kx�*�s�<��{�Q�ce	9�ɆEZ
7�I$`8a� ��������X
K܇B���Z覟�����G�	F\*U	�}`]d�ҏr�l@q�p�V�[yy�[j��K�'ϿA�1���T\b&!��U!����[���s�b�;F{w`��\�-���V.p���D�h�Wse���;�� ��ޥ�~6��8�Lo�����O�`3�K$��&��zW�+� I���9����w�����j��#�����k�"=n26�ཷ\��"f: ��^J�5C����Cgd�[ݷ��&�I=�����j����赤�]�7u������v�E|O���!T��뱽&���V*Ѝ�4�ZU��`_Ȗ������_�yO�1K�kf�y'��ZZ�PW��k.�O���s&Qv�J���R�>�Z[��ᇉ^�a�7�]�����ܦ���'\�E�w��=vGA,�	�>�q�G��o�-A��;��]���O���-\�$f{5xI�鰀1�`�0MZ +��J������	��Z
ʖ�ޢ(S�\�c�R�W��c:z
��~��6�v��]As~M79�u�"�֥��A�Ԯ9oP���G�Ǜ�貥�g'�&�{:
f}�#0kޡ��N�-������Ck�K	p�d��
��fλ�rw؁"���u��Xs2%��7��NF�k��O �������I�X�>��y�3o�#��+�0
�k7��y����?��D�F�}s�N�d�/f�?/s�G�e[��ݗ��%���j�>��1���Ȅ&>��*�ފκ��� ��<05ӄ!A�h@���&�a
����.�.s��d�]��e���Bs�}�i��b.������Y"=�"A�����a���0�w��Be��zj���O@��2��]`��B%���(�� �*7�{��1�'8���������E�Puq�^��寂��5�xf1\%~"�֓	�)j����O��ư�LL6{�3?g�|���D���Y^R1�di&���	$Gfm�k�S8dn����2x|m���)�i�P�ar>���/o<I���PG�$��ļ��c�c@+�BU���)��#¥�<G��K���R���6�[���!!׎NQ`��`�L�):���<��x|��T)51�"C�;�D!�����vAf4�8�5LG���&�BN���Y�x�2��p���A�Zr�	����﭂�ðCM�r,>�T�E<xEe�LY�V�!1KL�i!���8F��sz*�:�$X��r[�'�t��k��~��B�o?��}BL���~0s���b��X��D�9���6��G�0E�Td����Ǎ�tQv&꼱|9���u�1��l��&T��lwH,53FԪ�s��=�j/me��&��#-0"b�C�$�.���Z?h{�/L~cA����n��ٸq-?]�್�$`�KrϽ�_O�;a�A�����ӯ�}ym4���dϢ�Ru�2Ǣ S|7�c�h8_NFS���*԰L�b����Q��觫�� \���r+m6Rf���]�g�G���x��9�������Qi
_�6�6#�u�Yc�(C��%R����#Y{jA���M2J�X}������j�W���7ZQ4���a��%���/ч���	�-|:p��r���k^B��9�(�z"&����<���z<E��hfd�൉���P�y.1�`����x٢MyWW i6��4c�5��)�_�ݸZ�)���r����#Sq��{)���� b����"OH�v� �n�
A�<k�?������]ڔ��7*+�e�R@�M�?�R�c����:,��4#>)L!!SDz@�Bk����.*�)YQ�ZM=�4��m�[�o�G@�{TSs�̔@��Z��u/�x���e���Mc��{� �"�-�1����Q_br��"��xD��5���]�{����^���`-�c��̲��/��W�Q�7%B};+n-@|�3��7+l�k�v�jv ��'5$~�
mdN���1vh+�sv����pЗGQ��'�|�Ea��s�t�9�;>@�w�
y�ט_�SM�,��,��dXR