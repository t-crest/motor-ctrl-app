��/  ���O��B�	�LҀca�L�e5�
.�I����;�gʢ9ܭ,�_�l���c�pm��]��yz�Agap;Qܠ�]M���g��w��
�n�;0���+(�[m����G�%�:u��j�S�H�.��J���o1Ә`8kq�r��9�Y�B �I�^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK �fg�2�`��9M��柔nÓ�z��{���޳�#�����n�Ħ!���4KCǝ�0}��<8|��
����z�l
�a��@�:;�i7K�¿��Nd���%h��:����r�N�mI�gl@6|~��4�*����(tq��7�,ã����x�����!��ލ$�>���#In�m�T�d��vv�x��!љ�í�:�Lo�S��#j�'��Lg^e@��a,�:���V��d�P`,J��_v�HAx��+��]��q���٦qaypB�)u�e�k��;�j�~�JW�F#���í��G�a�ǝ@'��%"n~��7q�S��&�Lg���M����^�
X,NV�ۑ ;�)�g���`����W���oB>37)�>�Q�I�.�"B��3ER�3L���Ǧ��c?���zl#J�%���So����� e�gA'u�������OvN¼�S�뱪gh㴕;㩹��]�ډ������='E!:b����P/Q�����4�5P�L�[G��� ,'/[�k�C*�J]@9�m@�B]��٩�M�vmP�N��p��Y\�4����s�l���
�2�"����(��<E6��h���,Y�c�jL���p��}F�rw���A���nsI��`�Z�9����m�M�
'��6�X�*�!�ӆe�L������8o�(�8�N��ŠRd4��G�G���ĚG��x���
8�.���
��*_�\/8�� �g���9�W�5�4�3���HbY5dD��u�|���	�e�/|����f5Ȧ������ ���,t�<�ק!<���x�^���X���s��?r�ԋ�88����rP��Bw:�_D��b�����a�@@��:~�3&�h��d���$.���|�,�30�+hn�"9R��$I]��A#T�KU��')��%fI�:�NǰW���B�Pj{���D��Qv=(���LJa�b�v��~�Q	HL�d[�#7���:��1QeI���7.���qtb4I87�*�d�zA�BN?�a��񥺱4��1�Z��C����	J��*�Ċ؁�C}΋V�}��P���N����:� $��8��B4���[�
�FVi�C�1��0L�j��8����~v���G�������؁a>��R�V)0.�1.3���h5�Lp����K���_�Z���xȏnGa�E�3�ְ�
Z����m']�ǒ2o��̗��H�\S�w� 5��X�-���{���w�i}�z#~vU�.^�t�k^Tݶ_��#
|�̦-K�g$$%��G���@���e�J�<�i9�^�&o'��~I���
��φ�wڂj��W�����09�,�*��G�� s�/Sp�H�d5�\͌����E��ntq�&�LN�*�c:-�Zˋ0<����ct��-�I�o3��/N�O%?x�i��R<G��@�_g�˱`�1hn�b��%ikK�Nj���*?a,�6����(��'"�ܦ�4��)���	�Іj�0���4y�H*���n�o]h��z3�8�N?��+%�'������w]���nslK�{�n*l}"spK(J���F���lX:�1���N�]f�����pA<���خU�0,3��e�BEZ�<��#��i��0�}�r��\j�/K*�`k6+]o�Uʺ���J<<���吷V�N����ש�>��W�Zp2.���+��t#� n���6޲ڋO��+�}��q# �ݏ%�&���6�ɟơsSb�Z+|Hu`Jϳ%P��[m �0���h�:#��¼y�%�2��,i�=^��lώb��z��n��f���u�<��"ħ$P�b ��)$���ZN��[fM(fn!�\L4þ3WP��"?zr!��+��n�<�;�QlC�4R�7'|JH��K��u��fY��9I�#	�{H�%��h5'`
�X�0TS �@P����*���#���+�|�,�3�zK�[�|�!Z�q:B��y��T�M�7Ԡy����"ǧU@+�����䚺�=
��cu������Ӱ�7i+���M6�X("R��4�?��y��2�F� Vg�v����2���{���dcXd�6�R�[ 7qe, �6{%XOZ%�w���9�k�qb}@ ���b2Ѐ%u0�<&�θ�<��h���N�V��6��{c���l_d��	rșR��4�(Y�c��8@w`7�Ϣ�V�i���x���4̖Mw��"���h�n�?�e�fc�`�vLg�Z��i�A�+�%p�� G%����P���P��O����k1N��_2��V����=%��g��TL�1�)wT��R����[
a�����ڜ��k�.��n�~�����X�ƣA�Z�uKA�v8��bo����������� ���tijm������ˣ��^�#L-��?Rr=����W��f�r`^�	���V?���.K	��iJ
^�!�_X��zg�.?y������/E��`X�5�q�pۚS�	�t�08�1���qK ��g��^�Ɏ�>)o@Szz�w^h�`z:�8�;���y�XJ������Zү�p��0������hHe�g^aǰ�r�SA�������ɥ��]��3�Y��:�;|U���1|�~'CO݂#rs�(��	J;�Ez��3D������z�;7f_����7��w�FZs�=�k߽��C*(�;1�9U��X�vQzj*���ߥ�û�B�|9�q����5�3���#r��0V�%J�\� ���H�	�b��J�݉�D�?�M����̃G���<�2[��e!~���^��3r���J��{���B�L�������x�)���F��e�eqJ$T�`3[��BH��Ir�Z3+�h��a�F^:�l��FFr�~�ԋ�ͶI�2����]
�[@��BaŐp�ݶ�S����2�xJ����M�Iqs���܄���/��0��Fim�q�m���2(��i,(�����o��Q�o�hT|���9�i ��B��-�4�>뷍�����/Ҭ��q*��fŴ���� ���v	� �L����҈<���th͔�[i M�dˤ�Z{;��X���e��dt��5w���Op)_�s�ܒ)�+8=��A�jَ6��R+��ng�6B���č�4,�M���W ��5�,)t��	W� �:0q�?CtPlZ����f�s�@�h��L��ˣ��0��!�5����#��iP��;Cb{�ڃx�˜y�kIrLg����~"��*Y��N�Յ��ʩ�ߙ C�d����wC��q�2�w�s��z���#19����$����\tT�T��0�=�<K�!��v^��29K#��2�Y?>1�HG���ٺ����������W�H+kR(,��C�-�C���u�!��M�~F؟=�(:p����~�hJ���f.D�~e�u "�/̕a�c�1�ʕ"J��T�s�3��2^��F�D<��V��b�� ��w���^���Y/�W�������5ܓ �`��͜s9�֙/�ҕ M�����A�dT%�ce궆o��?�Q��ra�s�Kл���Ӏ��(�k-g�̀=���u��g�n�h@�[���5]�����/~�(�����ի�+T�����_b\�J�5�n����N��b{D9�����	�Y��P�^��s@F����0��r�k� ���D�'�����b�(|�i�%$��j�@V��s�h��Zy�}�ͲAP��wrr���;f���\�:��7��kSan��L�/�ޘ�b`+�P^��#k��௄�雙��w_�����f��s�����|Z�쵠Ġ3??��\|Ԍ10rL`E_K�}N���Q�������z�2���hAWo��M�ç!�W�y抈�
Tλ���׸]�ѻOX��5N��䍟$�)�֝�љ����7|"�3��1V�a���>gHΧ�s~�l#���-��ʟuoR�}-���� å����v��Qh����"�;Z"�S_�9�ؖ-vx��z��L�3?��&P�`5ˀ�eCI?U(�� S�>�96�C�i�ϙC2�����l���d��J��\u�u���i��R�����m���T��,�+��ޯ��xV�p^ '�2�t+D�0��4+��.W��}��=���Xd���Σ�C3��8�8�t��D�W%��a�ŕ��9ذ��'���GBOt_�V4�ھ��z!�j�r9Sz��D�֝Mi�����L����p�B��k��#����![�бnu��g�
�������������Qr&l��D]�����[/�'8��(D�o��<�с�r��C["Lwb)$�����-Q�K*
C�/��ƴѕø���mW݁������D܌�*� ����u��h�Av�
r9�-�Kms�p�L���Z���I�Qt�/��'���f	=|뷧�q�qR)&�x���E�q�Ge������x����v��8`�ޘ�ƽgh1A���g#�$����1Gٛ80�Vx���