��/  !f���<�bC]����	�H2q��@T�h_N��Uy��?�d��H�ؓN�F��)�
s�Ȓ�c܍���6\��4��p� �'��0�i��ͮ_5cd6(w�!�/�rb+��_:+��Q�[�*����CC;6S��k�;�N�Y|'�/��s\L8> �^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK ��3h})�e|���v�������� �M����� �(��_��U/�o��*�Mh��?�VB<���)xRb���q��ube� %���N(�o5]�%ۿV ���~9��l�K�!yD�#�;��v�T<r8o������g=���%�@/�]�P�e��KD��9�!c��f�~|	��q�=>�y"7t!QV&���]#�w ?!"�h	`)���ӳ��a����w�|ŗC�;� c���g�rB������ 3�vH7�oq_Ȗ�SY�\�)���?L�����`����4�SYF��	�g�J�`�Y�Nd�Ц��i50�+U�sçܣ��{*�7vSq8�HC5���Qfɲ��e�c��%PW=��r��0X,!H��Y�s	xm�y��a	\`�bر���:s:y�g�E�[��O�H?�Z�ϗ
k�����Q� m�Ƙ�T(��J2�RhsCDQ�ɬ���͐�}�#%xD��!u��,0q�����Y�����̰~'N����Sf)P��a�t��_�&�mތ����Ip)s���`g�Z\���A6���
�%��oG9M�6V�R=����������=;�91��,x��a%�/GEՀ��'&@\��{�'�JƂ�� {�3c7�������Fm `'�LEM���f�r���R��C��c(�;mB�	;`�Y@�4?�|@�:���Y^�2;��I�5�l\�F����əz��U��C�wM��+ɯp4���-^#փ9ޮ�r�qM��@_f�~�ݾKęnyխ`N��jR�&:��vo�>R,[�k�i�h,�ݭj�\\����e t�c1�ާ���JKT�C.�	nL�аz��o�>�1�G��D��h��!)S�c� X���t�\*�W�,���H�gp���!����h�u�%l<7���j����(a9�j�Յy���_����إ�� ����ӕ��"ٙe�i*u�ij9��3)غ6j>V@]�I,ilPLH�}�[��>���Q!�K��2�?��Cp�=��pS=r��g�$��[��Su�(��������u�%��������S]2��p8,��V&�� `π��&����N��B&� �p�n���UE�! 1�����1�;ʘ	��%'�M%6*���i1-fN���ש�Z(���<Ņ���՘���9-ˑ�Vn�p��쵀��o�X���$ ,}�(����%ϩ��S�g��<���X��\���]���S�i8w����� �F�3��`e���D�T�rj���\S�q ��:���D�l����U�&O�7��*��G>���YR�W`�T��u-,H�.�!��?r&����'�3��8��:��%e% �棖*���1��F�A6�M�����>�E��1�U�MJ�m׳��Ԝ�.|�[��r�D�X~�D{�Љ�XÄ��_Yf�}?q10Zy�1���������߱;�73�H{��Wk�Y���ɔ�_i2H�X���uz�9�ˮYl5f�N�ˏ�^����㡌H's�m�3ҹM�v<���3[\�����j�R=u�5�Kw,��9m�E�B�(�%�5Hꪭ�o�����c"�Ae!����I�{��=;�g�h��l`p����U�S{��S3J���U,��sT����6Q/��[r|($#�ލ�}��{
��ɩ�PP�sp�h���@���*�d�ֵcq���U\������J|�/lO����X�z��aF��w]>��#��2ů�����-��R�RPS���eI禍�+���U�u����?dA-��^e�ɥ��kJ�c1R��7N|�Y@Wy�F�Y07�_�Է�ͿD�n�ՐoIQ"*���M���8+j�O9���6���'>��H�ȯ���b�:�9Mr}�w՜��k9����~��/mk��>z2y����Lx|���=�,�
>j�C:�j	l��a��M�;}�Q��VS�k� ۦ�0c��#M[�C�� n�|�,)~)��z��Ṗ��Xc��W�hۮ]��Y���X�p�]���`�q���]�௲!kdflo�K��'D;»�6�B�,�FaҼ���gLf9nn�\���St�j�>�-V�9%M������><��� ��kݿ�~�[���{�6oߴ���_�7m]�?B�K�����ov*/�Ɏ%������;X��C�WfMJ��U	4u��7�8��fkU��Y���Y5��-}�n�P0�����E*`\Z��{�e!c�w�IM��Z6�")�����w������ g,�_��
;�bH�EhɽΚY>ᑛ�PJh�qMkÄ2&�F nś2��Dɯ���ħ.�z���O���$�A�C���x/xВ����F��Ph]2�4��6B{ F;2�f?��U\ue��YF�8޿��Vt��D��`�,����PTq�e{cKo`����{ҼZl��5��iݏ-��W�{�܌1�tr����[��S�?[�YC���bf}���j�Q����%�(�`���0�	�$w�V$d�
JX��|	<p1s�Аθ�������F#���b�r���.*R�<�:0i�K��fyY�~ �P��i��8�v'9���V�vY��ӱ.z��q�c��ytAjC0e�� X�'��������`Wγ� Ou��/��N�,���#�=��k\0d��s��+�S楸�g^*�j�N2&�/BW3�O�f���r-Y�9t�s�
f5��ƈ��{�J��:d[�Z��8��~TRI���V��G�9�h+���^��d�yC����
����ItC,�.�9�l���)/g=����|����P`�s�����D�)�e;ǀ����N8��Qe��퉫Ai��e����4Fy箕���Iv�@9j�X�z�]|���;�����o[UJJC�@�C�M2x����hµN�K԰�"-�j�72�F��fʣ� �k3���B{�%	gH�+�7)�O�|}��ǳ���?C�&&Y�����ΜFn�$Z�e՞�)q��s�0�n��&��$^r�mB1=�_��5[O�����HHK��ܲy�Ν�E3_�͑��]4x-;Vj�>����;1�N�ee�R���7zJ�NF��\��O	SJ>�;�l���$}�A*bBRqO'&��K��=����� 脸a&�}w�[�N�X�����|�1ɤ�?� ��������V/H ��!�
�W9���zߛ��u~��� f�((���t�f�r/Fh����]OΎ��	��z$/#������݅�ׁ=`^���,���m���j���#+c�j�M���1nK-�/'������rF���s��)-��e������
��,mxZSٸ4���o�Rq����I*A�g��No��x�/� �A��X|B��u�4|=V�P&/�[��_�
����Xt�Ԧ}"Q{u��Ak���cF�h��?!b�0���wQ��8�y�Z1�f��7"�O����#rM'pm��Éq=���/�oN�������'�W�r���"83.�۝+p7M����c����N�՘��Q��%nk8�K���j��׏*>c�.�r�Ğ��c�K�04�Ӝ[��[:ā,Aζ<��n��k�P��ni����<C%��Z9he"6�U�+H��,zy/���j��'�Z0��{�P��C�x�W�	�J6�52/id�6#c�yB��h���7�okT��p' AK[W' �~�,��^�_	W�>v\�]V��t�MGZ:��j�ki���W��[�B�"�A0[&2������I�y֞�:�S ˳�i��t��2�@�,��B�&	���}�6�����h�|��<�9�rC����sb���V�8T��TK7-��MSi���UH��sG]���"�/��s�.x�8�;��{)�: 
ܮ�Q�r���;�]VT������7~}/�� �'k��V�ʙ�r�A�%�Qכ�[G��ｘjH�$Ǭv8m�!��e��C�[
�ѬD��z6 �E�1�	c�bz����zj	5�p/&}"�%�
"�Z?��E��iv��a�{�Bqf�}��x(��H�M�ŝo�A{�F�5.��Y�#ﬦ�0���\�y����ӳ
3�����֣Cq〦��s�� ���WŘ��].� ����I&�J6����҇�~t��|���h�v�D�]`B-�7C��X���������O�.����w���1��\�X�[�O�,��Y�q����h���ם;3��D���I��bez)�L��t)y��E�[�n�<P���0l�X~���
f�w�`�sG
*5 ����`]+�F{!p�s~���ɕ�T�7��<����Z,���57�Rԛ ���F� �*�42�qO.�1��U��܈�������lR��U0���3�TkS*]0|]�����h�|�\q�(�A�Q�;�5�Y���	�R�h3^f��Y0�c���8iNJo�9%l=(��A�u�L��ŒW�Q��wkR����2SZ�T�C)O�3��?9�߹��S=��A��**Kf(�i�� �{�̞8� 6�m�Դ��*�?�x`eo���|0P��!{�
Qw?���x23�]+P��tz`4�(a 9Y.iէ5̞KH��?8={q�K�*$ࣹ�(�?�z�y�8��;�2��6~�sX�j��7$D�Z�)!���c��aX�cW%��A��OHM�[$lɊ��3��8	�i�-�Ӭ�~�W�Ϻ����4�i�w�:1a�C����@��!.J
����i%�b����)�,��`�U��I|�]U�]��j��+���+�N��(qC:tM_� .��}���<��+\D��}����q&��ծ�V���z�a�R�j8���Oi��D�._����$�ujS:�<���EiT�"t.j��y�C�яf�WuH�]�]r�%���>��+���,(�p���*b\��44� �E܁@�^t�+�m0�ɐ��UGz>�ύRǿ3;�CSdU��e^���&��+�'Qֿ�H���{������?&b�i35b�h���=f�L@#/p%>wb�]8M�ϓ���0ۍCD�q�k�F�����C�Eo5���s	�,r�Q�6��g��϶0eT�7�2�ai��o�̡�?���*�1�e�W0F���Y]�tw�)����x��?ݔ�[+&/�0�X,�b�,i�� 0
�
�x�I�3c]�'�T�n�4��gS��փ��H��.�K���)!#��VA.=���1���x�i̍��6e�	���Acd�"�I��0�b�C?��������DM���
�Dx:ǲ��
1l�+86c�X�Y�o<	��Û+^�p���Sb��}��'��qP���+�j�6�T�$����;,_K�6L��4ո�92��+�ӧ�� ����S]������kc�G�0I�O9מX]�]�%� 2�ʸ�1Ns� mc�洼\��7���n�Z�/�bo�T2I�5���V@��-oz�}.7�9
?�X?t�}�b�1�a�*#�&���^V��{�gn� ��B�X�y�3��E =���?���P��'�2Q{A�r�]H�h�1���S�;F7���~h#��G�λs��`�sXo1���G�`��FL�EA*S*�=j�*;�lvD����� �+�m�q�Z,Ψ(�o�%��G&1D@�\�ʓ���ѭ5պn6��&����� �1�P�RR�Ә^����t�O�^��v7����u��:�G�ǫ�,��ܓ�g��!f����%��ǎ�SI�	�R��,�=�`���������i<b�S,X�� m$ �'ړQ_�+7��	LT�ei*�Qmp&J.��������lI�p��x�`�/�oC�o[��| �V��&���l�8�M��n��!�Hezޏ��a�DBw�d݀ǡ[a�Ԣ�P�YAnAF��dJ�Q�2`я��	�W�"C�Q+���$_�L�얓 c��i8�RW�<�w���:nL��̤4K�4L�x�D k�
쾗 $JKLl^�M�2g�7b(��ט/6x�9�틞xhh^��(�j��;�	wU���XF%BVc!�>�����i0V��@���l�}�'�:�N"�x��b�5�ŵ9k�_`�9�T�'/�;�4.�?ctLX��ӳ� |>�p��a��`a��I�R	��v��R���p�^˯�nY���ЄO�w�� �Wv�ѳ�nUD����O��a��,������o���n$+�<��@^��8�ؑ���Y<�B��s�ߛ�:R�ޓ��>�r��9��v��%��qEK�GF�l��#�����8�'���^}�?�|��~����\�w��1��C*��eΘdd4�<7hV7i8�`�mmZh4(�U��+��:�E �m��:+��y���aP2��P ������R��sׄ�)�����9v^�͞'��������H.i
o�v�Ϊ>B�Qᡫ-B��&��5C�>�/��=^zc�N�G�����˔�r �cW�D��O�>�x������_{S⌎���W�M�ݞd~+�ݝ�b2�4�A
*���Y�7�||��1�F��h&F�:-0��a�m�%��^"�"=ő &��h&�����	���?��K=�	��?��a�VH���Y�$<�K�yq(Ko}`ose�dO�^34Qf�ړp�� �L�CA:(��9o�=�=q�=��$�� �4&�@'�~���AOO�v65F�`�\�����=�F�0sz��Ŏ�sY�b��I5J��(����1׿%L��:��@������9R�`�fݸTy\���k{\�념�u�sC���k9��2��L�� 7>���մ,�k� �A�)�~^+��O�����Q��hfG�=K��tW�[���wJe�6�Nˍql.[  oq�Y?gڱ�j0��0�*VH�Z��+;���	a�`��Z�[H֩�L���÷2T�|��AH�l�Kͣ}�t�������+׈���Xml�ڝ̚��܂�le�%��#5�z���j�[P+�T�*���g��<�n�y����Z�Am}�0'���'ö�[���7�ˊS�it	����C;d��y6�@��w�Smk�[c����EWS��*R�W��!��x(����-�TH������҅AҬ˞0Lay(��hɋ8}���'�(T|�c=	.���r'y1����{VF�5��[�J�p�4kڕ��c_X�D���|�zӤ��g�cEM��j��p��i�eΧcM�C���[`o0c'w�&�A���A���l튪��*�5l�yݒ��-P?j�D ����P��QlT�9�+5<:�jQTHr�ْ���r������m\��]�e�'|���Y��-�;c����K��QA`�������:���J�՝��B�l��m5i���74��P��1.yp;�LQ�{�OC�����E�9��K@�-zϝ+w"|Z�p��;2CC�T�^�u �aH,i����>�;$׾���E-�jf9��ٍ�۶<��.K�m��$��j�G��z[��g����Ý����7�7��3�͑����#[�����9�v��R	*�2��b-s�b�g98 �pp;5�Fɯ�6�/$3/���y���}���g	�(�de� ��Ԑ�!�Y�`��x�Ӈ�� �9�]}R�v��E��>bN������<�N��Wc�QÒ5ѤW�k7~ڹ��'i�9Y�&h��z.�r�����/��6��/>�ȷt�ˉ�**�uf���A���W5!)?����!j�v��喥�M����XSAB���z��6�BU����Rʳ�[bb-[�X&#-�K�)� e��Ds��f��J_� �M�HP�`�����1G�4\do��0˾�BG�F�G@j�>%^)ц�W�U��u�O��i��t��rz���5)�C���!�H��m�]4����ڒߕފ�K؇��g))�O�`FF�V�& �5�OW��#aE���44mF��1��ۚ�HZb?�_��hzTL!�V!��P�"B����LW?!@����
���)���2��-��fy�f��\9�MQ����o��A��~]����'ߴ>
D�Z!�>[�u��g=廑v�"ȍ��;��_vW[*�d��	#=�	eY=q$�=�oc~�z���w��yI�/.�M�`��3Y�]ȣ��7��>�+���@ۅ��Q��hV�g�	�b�_�Q��:$�{�K]���R�1��斄O3������`�����'F�e�':Q��^"��עa	~����x���h�zY��Cl~����qB�?ߒ�/#�o�&1�}~:�H��5;�ݥF��|��ޛ�0}5kbJ�tc�?ģ0$���S�E�@�V�BJw3c��jwǜS�.S��͗N����f�9*􋱚��z�3|%js���q��J���x'��poCǯb3����R�r�W�W�gK2�jm���P����\�;:ȱ�[������_������|��}TVP����1ǄnM�����t�b�����e/���JS~͌��o,J.��UC�Z�V����B~[2R��;;�hq��c�̺y�_�C��fB�'�e~V6��x'޲&y���~i�;���"������R��X�I�������ׁ�����Yp�f�ܴEl*�����>����4qY����6�8#�#�>ٸCE��q�(6�i�|l}�p
f�.n�2��4�u��wJ�O�:ƀ���cW�2zb��;%���l��2b^��T� ��e�_�v��������1|�����l��Ǵ��"��r�J|�:�����?����m���(r�r����O�M
�
�g�U�Ϳ�p��N�;W��.���W�����3����_ �؀�R�>RFX��I���w��=NN���=�ɢl��}�Gؔ��2E|Mbiő���'AR�V��"n��R��[������M��ˮ��	��t& ���?6�sI�?v!;���ru�~��cf@��S��xUXׯI~P���}�^��Hc¾zʫ���0������d����g��
�!H�+{��e���T:�v���A�N�+�=8��5:Z���(�c����#�]���F�l����#"���t�e����h�xE8�;4q��@��8�ҰMXm���G��vيH�������
b�{]�'�)��09��ݰj��:�j��O=:��O�Q�v{�d9�}ۃ�2�b��L��ٿ,I���I����g����p"{�]�We��\����ݍ�u�!I�{3�QH?(AK+D�~~���&'�욘���&���?��Ϧ�X�	G�eR�t�uf����2⩍��6/����Xa۩���l���6՟�~�������:C����k�:� o	��.���1)��\�-��6y�ۀ���ł\�E%�rX�;ߗi�"<1���m���g8���7_kA��5ck���y�+]t��y���;��6*��wţ�������0��ՈJ�I�����Fv"�HK�V�2��?S]���]3$�U�{ٶO�kCX����tSa��/�K��{�p���kJ���kA���+��0�]�6��篨�p�/�pq����	,�N�p�K<	ҽ���k")�<��HT�^M�#zҖ��qn����CH��bpx�=�dH�.N\L��~����g�nYb�}�۟H����m�]��H�[�z�K�,i�����Ec��OUMQ֍���2ɸR���jA��؜���]�!\�P�ߚ��k�ȪN�~�u��Y�iu.�\��{� ��В��׹݃l��Jh�5G�w��\�8�MS���Ꙗ�i������FC��d�
,蟡"�8n>9�ޝ�i���a��HZ�M��G�a�H14�mW[�	"��
�]QH^���ΖΧE9!�̲���-�p�J�q��o��Ͳ��1}N"��纨T[M��^Qot�, �b�2�r�P�"pm��N��OF�_O6��s��\X���wp��pUI%/9>K�[�o���d;P 5S� �06�3�+�-�QV8�SKJ��KA��Y v�"� ��٠���BP4j�b��`�{j���J�(�[�e�@#hP�l�Nx�*_� 5���&O�D�tO�)�b���H���S�L�^�c��pI�|�f��#������j�/)��d-�J���E�%�|���+�����̲�g�{��	K����)Ӡ:��󱳗F W�B +�J�AqUb�d4����/�mQ�g�ڥ*?��79�P�]4�V�����oF����qv�l���b��v����Z
��H�����GS���5���}=*]�)<Q�%+
�~w&g����p��
�!O���b�����9�!o�;¥��	��,1��Mh�D�fVR�Ĝ�'N��=#}�y��@�-a5`J�hA&����D�y�f�S1=S�"M��@����W}������ v1��ٕ_5��s����Y`{�i��}�:.�<t=�A��N0R��_�yK%~`�nNC�:
c���<<V~�5�.�P��g���hK��BoҠWɠH�s%;�m���k������c�#0q��X/ ��	�r*��RO�.XQ�G��	����/���V�	:���v�
��WH��#8Oj�_�$"}�� 9y�ܠ���F�t�y��9�����;�2�x���x@u �7�3s�խ��@���	Z��k�;k��Z�<)������Ɖ�BP��������F�� �V�m�����	�A]�W.K`���T�w�ET_����6p~8	J�%�@w�I���>�*o�q^L��B��<�?�D@���#ԥ��v�zp�G4 �a�XcDŷ�'N&��4���I�1�6�:
n��jw�+Ⱥ"z #��#�ǣ���ۂ�:�"tQ蚜��� Ѩ� F��+�֞�t|�����a�)V�YY:2+�OE�u��?6VJ�?�oP�lʝ &1L�҅��H~�|�K����^�:����"mA��4�K"WkS�g���� m�h�dK]Jk�^��A��7M��;\�X�m��'��G�&vy����q2n\vO\�<I�N�l���y�����Z6���(�V�h���|H_�л��Ì�w�M�a��k?Vv�n�Dy���d�����X������3��~|"�w��WN���Y|A8Iu��.^H8�
�1��LFFU������^� 55�Q�>�Zĵ����O]MhoY�z~����w���PR�k#5�͗&�o^����W�,��]e�EUo��d��wI���0/;����<��Ҽb5�����NLl"�<2��8y�L�t?�e�
���mc` !��c�?�x�͌�����E�:�Qi�#��?��J�]�	�=�_r���x���>�1�A��#�#r(�*������Ќ 8�-ĭ8�v�NHZj�q>Ѝa|yFt*�O�dv�/!Ӯ�$N�z;��%�A�W��¯�u�8��h���+:�Ѥ?T#?ܚ(���4�� ��ע����y���<�ĉ�L9,C7���)�]u>5��:�R��	��H̖�58�W��} �S�G���#3i@�0�������Z)�!l*_ew�MuhU��B�������"D؇FːY�e�Go���o��0�o[��j��=����z0=sUGHh����J�Y��}ϰ��e&wI��+�����5�6b�c�G
�LDĚ��DY��ެڷ9�4gb�Ji�o7�6�����ݘ���zA#�ؓ��vLg4Q��_�P{5k����^6^A<<��Ga�-^�w��F��|W���U��|�mf�=+J��g3\>��7���ւxY���9�)��X	�ҿ#�"wt���qV�>�x���|~֨�=��C�h&��JA�Jt k	J[�]�`$���͹#�a�\{�֔�[^����Ħ��W���N�&[�>��.���k��8�"�a��-�z|)A�N�=�\.~����Cw]�}�y-X@;$���'6�K���
-d�q`[�%L��y�ωO!z+�W��%J���i�gatքѹR@�R�JZ}����p2��8f�%6c�K���M��ln*�zG+��P��H��HT*N�tU�D��ь���{D��7�"�o�S�U3x����%[��7҇�yH�h	P��,���6}?}��f6~��2g9��"��^��cR��녾�ɜ��$�@��4*�q��-���C�}2���k<��G�E�ʑ�.9R2��#�.��T��Z+�U�"�榷Ñ��1�i�c���� [n���D�F�C��\+���9�ݨ̏��>,] ��kr�E�Mm������3�K����Vf���8�
����!�M�s�(�:r�]��1�끦7Q����Q�4^g���9[�;��o魄G.z�-��DI�]�Ň1�i{��F/����o%JL�.��t#��"u�׌�|k�t
�*�we}�2(���H�*�aKH�S�Y��C(SP����2�Mz/� yD.�~>���Y��(��ŔI�`4H��u�RaV��b^���6���e���,����	r!^�G���}����Ap(�.�9^79�-Ova��v<���3��8��zh�Pv3j��G2���ǟ����}����V��tf�/(`�2�BX�U�3��^�k-�r��$�7��46A�ih[����מ,�C����({l�-�?<q�I����v{�
ܧ�}PO�6j0=�V�a�$샙�O�q'�������X�y�]��n�nYS�?#�l/v~&Bh׋q���?͜j������og���6��}oߙ�LP�I��:d�c���È���M�c�Q�VP�%9W��C�σ��n���70�������~m9r�T�lO,�-&��u�6s�JDG�p�V��_�ye�vqΝι�S[���Zi���Vd�ꞐL+��ܦq2�4c���Y�v㿑c<�"z�Y��s�i]؉�s̘ѵ��"M�R��\�(�g���-bE��lD�(W��?�U�]1�X��a����0�h��������b���d\�&�Ć��]���!�S_��d2hҴ��J����tR�E����b��8{�q������9)�	9��v�專|-��hD\;�>�|��\�)� �����EK��JK�۲�!P�ѩP�죝q��R9���.��cWv�xst��y�֪?|-��6�"}Y$�$Т�J[��K�U��=����=X�6�%���x�,S�z5���v����N�l��ָQ�����`�9���K�bK�E'}� nʕz��Ի���酫$�9�B����I�4�W������7�H\`z�vF��e2�ܯ�PEa2���Ci�����z��(��978F�`{��(F6�����v]�,w���u��c�3^�|�\�t���ո{�?��(�+��G..�=�'DcKKB7m�铓��4w(o31ēƲ�J�W��4�f,۸�9�$)rZ���1�5#�P�&n���?�SҼ�E\��{bn`N| ��p����S_��'�}C����u"0B�K�ô��vH�P�V�f`}ju����<�M����$�Dm}�݇t��	���_�����:u��x׼���Y��t�-�P��Dd�@-@���.ml�Ӝz�6`����n���&9,��2�}am��ه*j*cy���׻K&�3�O";�=g���.l���9��_WE$3�c����=[�2�K���i�{H��/�5k�����K�ֹl�F2��&a�a�$�L�+¢��p���`~t9�E��k�*���[ui�-o�܊۟3C�����GJR����b_!�천�ED�Y�DF`"��O"B&!Q�Z��iG�D@G�
Da�zj�-"�S^]�)����z3��(6ڃį��P
��������3�;{�z�
�K:�Ǽ�5,v:�i�dE]�tt(u��ǹc�Y��H�9���X �cO�ޭ��L����L�#��@�'��Nղ����?��/��o��ԯ�7) IIT`�UV1� ��A�4{�wX�7۝�|��[HҬ�%U�>�� ��|�N��0S)�d��f�aY�!�FK�c�X��m�F�z��N���g��w4��u�Rߑ�Y�%���d��C�T�W����E.����gJ*Wm_o>����#�T��\>��"�~!��X'fG�$f�O�+��#$�+$�*K~鬉eJl6�B�3��dg��ƥ�!b��Nܭ������m���OH}��@�.�7qH���S�#|�w��N��~�d��m>�p��XP��8L�5���6p�d���VKSV?�w@o����I{i��I%5�~x�/� ��x�6��gE�f[�$'�T�ߩfȝ����E.�z��;�%���%���t1���?��)�xW2��>d��%���Lq1��d�|�i5�'��Eg<7�t�ÎX�M�d��ӫ�����KxjV����,4�}4�p�-l����}C* L�ي5�5�E�W��꺌�MZv�k��]��L񘓔��N��voy�j���L^6N:�)1f�r��^�cL�,�d��ɤ��5U�W`-����фE4��b+�@��"
t�m件�ilW��'̠�7Kh������U3���i�?�] ��f���Z�+j!��L��~3L�GN�-�x!
�R�r�kF���vp�z5s�"��V�֯a�\r颜��-��x��+uŽE���E<�V�"h=q�B:���b5�tF(��гA�P����Z�� �B� �^at�E37�W�k��P���S�|�k�ϛ��dX$��;��qn�OF�4K0�d��9tB���
���S�HOh�<��t:�ʾ��*�ll�O��b%7�<G٦s�
�c�(&K��{J��ߍ:l�ʄ#��)���+��$�R�~у��0��Z���~G�;�O����$�Ė/o�ނ��r��1q)	Ș�\��¤ �=E	a�t�*t#"��Q @�l;%���(�Sq�Y�l>�՘�z��oX��g���1;�{dV�D��<ƕ%��]�r9}�t˸�o:K������0{�S�)�8�ѕ¦*q�-�;�i��*���q�.��T+���Q��[
F��� �&��1ĩP\�2>�nA0����@�ȉ�����y����)M(3�a��tr�����9��̂�I0А�њz�PC�{���!��e�5Xx8+r�Y��N%:����Y�������H ��i�ff�%�zXC'��$�c��~IJ�i�a\��n�}�H&42ZZ	y	�^�k�Mzf�j����n*�����<(la�&�5x;� �ㄸ���Ov��Q>���s�N�U����՘�gU�J����HA��"Cyy�7~,.���h*��Z	 fʀgԋd<-� Rma�b%y��(q14�Ko�*��i;���b���ֶL�q'ś��-J��;z>�L�|JpO���0K@ɸ�
�9�v�U4h���$,�&jh����g�"X6{m���Qp�?X_�����:{s5�$粝����ұ2(�(�G�'��`n3�@�Ew��1]�ؾv�1=��/Fo���<AN;a�=�D�����2�n�&��y \6���uo�ny,IDWz��jU�����ZٍO����L��./�<�)4 �K��l2������7aUݲ�
j�tT6� ԅ������F�M��	-���b�,��)�:����	g���?|i��~�a ��+��Q�K���_i�P^�]��:�y�&I��%3�"��J�=�Ŀl��g��g�l��e�]�㇤O�MM:��^fu�M�mkQd�.����%f`j��o��l�Î�=�"Μ'ӈ[ �Gt��o�r1�q��x�?�^���cV0e��2q(&�<��"���= j=xD��K�K�'�ҷNg�UH��j@�Z��L���b���NΥw�C)����R���+rHhH!Ӄc�hڗ	���tZF��n�JLWCv���(�|�"��x��_�#�l��w v�?l:�,�'^Q���
I��Mz��.����ǰwů`j04;T�����V{���/����]��z�6��-*��/S�pWU�Dn� ��]Ʀ
t� �BK8��Ս9t�No��ŏ:*�௴��Va�k���S��Ggɛ;�nF�����v��Za��0�,?2P�n���+���ost�y��;�~[��1��Jl�S9���=� �'�hu0��tGy�>JӃ������T#���k�n��ˆ)Am/���M� +�?�7��{�F�iGw��xI.��V}z���c~3��l�+'Q��.h���I�dsRLeb�a��3�9���ق�i�7[�]��d����):=���#Z;���-M}��&�H1�w����N�@:L(+1�_��(*]�'t���?t�x]f���f-���^���\`�k���m���u�!D�1+�V� �GCͰ+9��X{�<o�IHǜ�b`x�Wt<LV���j ��dz
y�uS����Nt�&?�u�r{N]��~*Y�+�MΫ�]&�����3$�I�G��1}�]XY�3Y�t�[.��������Vϧ�X4w�����7ړ��@�����I0��:�}���T�
c��R��|H�H.�q��<���)�b���S -պ1#����o���Q��)h�_͘���1�0�Jv�a��3�!�h�+�s.i�{c����g�)m�<'�I��>tF��!9���r�Yg��e�6� *'>�k�f��AӚ�U�)�L�B1�ʺ�B�<r�!�:�[�øɢ�&�8A�������<��7�T�m,���k��ݥG�&}��ؖ{"X�g����Xw/���͎�|Y}h?��4�=�}����j%D�;�=4��/��	���ise?�Jt���8��ә��ӻ�D��4��o#�S�%˼�����zaĀ��M�]̈��x�kT�#[kŎ2�@��7�4c�o�|��w���i����a�K�����Q`G�0 ����Ñ&���w���Z���Z*��y<�l�g��\{:��@���8ٶ�Qo
��E��ܒ���ܝ�g�gٽ�3� B�V`��AΔ�p�'� ��X�	CTS�_zMl몂keq&�\~�dNvD2����?�,�ٍb����|o�7373�D��
��_���2���1	��F��1��1|3��C=u ֪Y4�M���É�-[�q\�Dt;��������N`�f�~�)��у?k"}Bq�rz��Q��r�F8�D���4���*�d<_n
�iSC�T�L�����n�5�m,�I�0�#�e�2\E�M�.�T��Ѱ���-]�{�=+(0p�o�&