��/  =z/m���z?s>?5��B&KN6:mJ��B�\w�:B�����g.b��/�XJ�;�P2�6�#�Nnھ!��|�kǬqy��"��#潀��)󖻜�ob�,V�H�6]�D�c�6��b���¥��.3e�0��6��;̆;�b�;��AᡐK>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�cǖ�x
�Ą��8P:`�((�w���岖�E��
���Y��?!J���j}�i��a�URBҒqT���fW���M����BB�:u{�� 6��oB�;������#EV����P�O$N���m����t5ckƫ�n�n ��I�ҾK�*���d��v�����"���g�o�
!��g��y��֙�ˮ�-����w�߭�SYj_��˔|��2.dP�]|�<�l}� ��Q���hA��5uĭ�%ʈ���-�\�,���d��M����h0�������6���7���ؽ�'���x���6�.N���A�~_&c{O
��t,
Hc�#���1r��e:V#���K�Z�^�N�T#���Za��	+?��QE���Mw�5J;+>��I�R.w�\���(�x�ё�x}�����qQ�p�Cy�0�*wN�˦<b�I ���8Z�͇��I�+���{nh��{�ncs�(�n��ǳ@軲X��`�Aߘ�GpX�;<�����
	�7y�	!{}Uں���V��F�w�G�rn �(�wOD!��^��^2�F9��N�K�㍨�������Х��W|�n�}�ҽ�UD��0T����<a5IU���/����j�,!l������� �)�meP+ph�J��5��;� ��〥�-iG��y�m�':������-�S#^A���H
L*�T��uWjb��Џ��8�Ob���wu�
*p*W[�{ůX��{��y<^Jpx���C��5���I4GT�Mx�XƖ
���0إX����Tb ��1{���3w��;7d%~�+Á�Ej���ͱ��D'��I��O��ǒY�F�FTP��W�W	��LX�핋�ҧ�<�;~	�<�\�e�����K�avvm���q�dX�5(��*����� �n�@ؚ�­�^�p@��g��IK,����3�������:ݙ�Ǉ ���~���6x��-!J�/��L�����!::�q���ERj7b(�r�Ͼ5���J����<�ET�҆�2g}3�~�������XZm{0�a��p�7��8�:�f���(B���LA�_ Q}�T�B��I�oY:0���b"�3`ߚE��<s#Y�qlm��ѐh��b5{���gK�4�n���E(��{41��8��=�v1�T|��|0Q @�F��r�я���=3�>�M.��8�D|�&@`a�~]�U�����v}f9����0��?C[���b���4��5څ>�u���ҿ�ށ��""�%�+,��ܻ��{Qt\��'�@�)�D��z��2j��^�4��B�\kZu2�F��^���%�ɷB��ɥa�eu ��� G�L�ى_����fͼ{#���5ڥ��EL���E	d"�^���� �A۾��G%r�7��j?��PB�����+��oB�i0�=��-�ŧ����S��@8�*_n�FT�O���!�F������{F����dS���۳�ECڮ���mw6�~-�gw��8JO���R㝕9HZ4B�Y�����Zb��o�4�����$�Ē��iw��o)��H0��8�%z�	����_J���{�iQ/9wwT�D9�ه�����E��Ѐ�[)���L�W����YUez[o����{B(u�~Ra��w>���2Ԯ�1�x 1J��C�q��m|�z{�l�l�Z�Da1G�b�2����Z�5�_�D�{����xYi�Լm79i�����d�`����[u^���q>Jn�	�'����^�h�i�By�mSy�S� ���K(=4�^�W�.θ�~Z��8J��� �\�Ė��kCh~�w��B��>�;Er�W��q���^È��R��lT�\l't�$���nfz��6c~�{uKT��f�2�>	!�֩���ǚ/���E�Ӹ?�wӠ���3��+��n��4��5��̎�X��u����xP�%~B��ŉwǬ����Gj�W�����p�w��u 'N�u_F��}���H4cTD�d4�.�Yl�OF�l�>�$�z����SMMa4$W��3ƿ������8�Je�٤�o��x�{�9]�W�ψ�B��4�]�Z��J����&�U��p������a��}�v8*�fC7�D�%l�W����do���OD�_%?������KPpR ����ȡ��;��{4�$�N��
�>U::�0��.��˅
u��.-���9��Y�5XzOf��p9�����_p14�N��/�$��%���W�150�p�u{}�W�0��t���f��S��@j�ʺf�F��4��d
��(������w��>�Ҟn��ę#�A�H�),ӚN�UI8�J_�[��8�Tӳ�ѯ�����ի�9�Moli����},6 �#�@,b���}��1ն�+̥�(9�s�*u���V�4"���=����F�ݐFa\z���	���ƿv��z'����!�����~���/���ը�K�J5u���=qҸ������K�J�mP��a�-ߪ�/y-��4#��>.r×�>h�'@�ue�54g:EU�=����(��sΣW� f����$��b�92=.��`�����?X��VL�ѤS+��$�G�.�n��vM����Q�]�P��.o"��zU�����|��
�#�'ԓ)gڒ��?�j��g�e@�^�O����3�&�,�'	�e:���cg/�t��r��a0����e׵����Y���/ݙ���E�sb��-IL	�xܙ7�=@�Fĝϩ���������9���8��U�N�UY"�4K�2����*1�t���q�w�Ã��]��!;o���s��������&J��	�x�y���`�s��dL5��1[:R�3��W2��'a���#���=�y���>�&����Ir��zit@�Ywh�ӎj4�<�x��D0�oiW��3�	m|v i����xZ�d�.YI.���U�2����+�#s��cq�\l���]����B��z2�����fN����M�>*3��E�c_q��M;�OÕrܦߛkfU��&H<���N7�ZMI�+y�Ґ#s]*�,.�G'`~�r ������S�x�>&A�n@w�#���''I� @M58X�^*N�,u2�gp�t����*�1>+)	cE�텟(��&��%�t:V(M�z#H�4� ��N��ǰ�17M,�,�|��F���NK��
/sW����ftL���a�&�ԇ��_��+(ʐ����`n�6�b�9Gi��|4Om�F�bEެ�qdiCtD��%7�^��u���}�m�k� �"��`>MP�|n�;.�Xv����"���M�	���A�'#���q�F�X�㶧T�RR�C���!�?1uV�3¾�gxh�I:��Vjy�2�V��r+!��c����g;��ú��+t��"��dY��;|��629Ì�rg�"�������G�R3�iT�gn�ơ�<@��p�z?���+��2�i��5x����*���5��Җ!.~�Μ��?iq/ؔ����eHi��\��[�~���ۍ�rؼl~�+(�B��˧�"�n��1O�NS�I�u�e�Nx���aE�����ɺ���eJ\.�Z˻4	��gqPA� ���D
�c��ı�gj����V��߈�W!���JiE=NRR���@���w��l �^A��g@��%��9���]�J�Wgq�9�>�v.�|8){�Y�h��W2���yڦ��	��!�r_50Y������H�]�wYbЧ8i��L ��;�"��~1�/�Y��XqbØcl��b$�DfhὡvXi��kͮ���RJ����7��p��e�~�K������ҋ�;�"��
5 �4�-���Z���ީjW�{��^/̡�9t��J�RG\�(Ư շ0;���A�۹�1^<�K>�C1���zp��ya�����=PS�N��"�OW<� iI�؂,�-[����E�~j��W�)�Au-1x���JT"����{�'��;I綕��_���1��(��G�,�+g�I���O�~��WL����A� �/���Ͷ.��OJͬ�@g��Ep��e(�R���3����d
*6�T����yq���ڞlz���L���ԡ�n��LP��$>/�bj'��<��+6�r,�̷O����8��\�砚MZ@�P�9�!�n���������VpI��z�.+�N���j#���d�Dc�`v��Ƚ>P9ֵ�p�sȯg	r6W��*�q�WL�B�z��k|��DB�)���HbV�]��o/��n�`�U�Q=�1���T��ݬ��&��},�3�c~�D��k]�7�rc}/�Z�Q3��i�D��wr�AĊh�|��t�Xy�r� /�Џ{�x�MGr�o���PJ��I �b �=9S�C���Ui�G.��T-�[R"`���u��	�1����Ƈ�f�ߊ�R+l��H|-�%
mJ�[+cΚ���I�Q�ͺ8���M����Ftϴ�O@�n/f^5f�ɕ����_~�#y!���W:e�9�Cwvcb�:!�'V[�qU��uL=�c)������[r����9L ��IP��(,#�lSf:�+����mv�(�~i�p��0�?Q����li����	df����f�'��ʸ�ݶY�7��z0��ߋ�ص�	U��g�[Q�����B�;���e)0	�'w~Ee�e6L0���(��f�"�������	��+���MjK����jm�����0�5��'�a���_���>����#$�$��wZ�kI��Ӝ?��V:a������9�9i�j�0��-ڊwI�|���wٚ�����F��f�3��
�m\�īsW#Y�^�@�ӵģϺ��	��	�1�D]���TLl��D���k
m\0G�/�ep�3p+�/Ғi�5|�Z�il�^r����cZ��k���D��-��kڽ-�����)+w[����C��L��ȷ\��s�� �\I6vr��p[!�����.[�Y�x��W+�|��#���%�ߩ;���?в���n��&I�Wi4�Y'73;�����(r*��u�&��h�ׇ��[��x�~�9z��v����ꈜc*U�Y���-%m�g���3ϋ�	\�4)l8����L������9�y6rp@{$8a��@ե�^jaB�.~o���R@�!Lg�~��gO�pع� ������B���5�JTq�ǃ�h49���k�f�.E%|� ���D���|=>��N�	�0�G�Y�I�oΤ�,<�X�bM�����ECvF��SjG�n�M-D�t6��z�s�D���{�o�E+�=��2�&@S�G(p_��|/̨~�(I�@b�ʹ����|=��BXj�]);�}�Y��E�z��p_��,��ԧ��t+����`;�6�vS�Ӭ��	�Y��`�G<u�t�N@�}S�Ϭ��ɵ�U9	��
��3AG2-%��F���3 ��1�󣘩��J���v�g���Bk'F�cp�2j���L�v{!���)Z�P�uD��~#�)Y���ń��M_��f���9y�
D��H �P�����a�����_Y�ݹ������eF㕟)ű�ǖ*>�N(���K���=R�K:4��Hu��"|w~�;�f�>���T��� �=?�F���Ŏ��3�Z�5��(	�bJ������Ǩ����.������p�Z�|��9i�
D����5�s����(9�X̚��߀W5�.6��u>�O����S�h�X��!����Q	���^A~?��Z��X�ή������A�1n�����;"i�o�n�(���K%S�5&Ċ���V���
���0y������B�?s+e�g���W�L�U'�K�*ѓ���b�c�	ݜa�>�v?|l�gPr�\_�>��v Y}1M���Lm�_qhw
��O�O[ ��j�y�5,�q4I$�3�iu�t܇��j3�P �!�ӊ�n�d�{;y}�DP�ڣE�y�2����4q`"QQ�9��9#�c��ؘ�<��l�"����g��cp�xB�����ϫ�q���V����ŭ��v�o��z�t�4z^�u�`@�E�G�Wa)�D���w�5��3�9֠x��t��V9���[6U���Z�]���g�ޝ��u��ٮ�V�����~�|.��<��Ϛ�|�:N�٧'J����PL�
:�ʩ%����C�7߱�rog�-�g&��b	 �N��9�*8z����]�FS�K�؝5Fg���g���-9�l*��^�PKE��5����x�O���J�C�*��ZC9*aV�U�YFִ��T�:�Fu�<E�8����z��YA��r���Ԝ�[r��K=�B4͵�����K��v�im���C�C��U�EJ4�>Rv���7���2��O|U�_�>ԏU�_�&"��<�p�Ъ��q�B�&��r�X�`rp��;✆(���
�����!��S��q8���Ԧ��E@���@ގJQ�%K�bݼ��e�G�j�15�#2����/��d���G���^6wbn��`����'�1�+���|a1a ��#�m���=~�f�X�d���f-��G���3��g4q��1r�=�N�|��y�"���F����"������P��K�T@�$T��Qv��8��-�#u͊��|[5u�8g�����H�x�!�`*���G��&�P��q� ����_��P1���E�.~��Q���1��9�w�}e��_}�l8��e�L��7�;�X2TA�����x��k���yH�G	~���cú=���
��a�B�N��1�j����1qf�2M���%}�^f>���M�r�gO���J�RL�t�Q�������c��J����/u��b��1wD�̸�P��'lͳ�O�27wB��k���p��R�sM��-�zߊ���֓�P���WJ=�[��c	e��,�byB���A����e����L6��,{ܹq����?Ag�
œ�O`VR&r=����u��{�;�J��'W�p�\�O1��@^+�R��,۟�u���b���es�0F3X��	R�w��᭶1��������;�+ĳ�139��":k,2�ѯr@�LQ���ݤ:��=�b�ȩav��KS o�L�f �}�2�����EQ2��U o��Ǵ�Й_H�w�P��\�Bkf�(@�g9"�/�Dn"��C��_5�<�6�T���u��zv�/��(�Ë�qT�>�!"�"�b�*ꑌ[� �����UTG��%��6@,��!��EM�����~
�v���ΰ ��h��|a����J��/(�R��~�U�����Q��L߲�=k�L�$����B�9���4Q�_��pACT�Ё>��Ն�"��4���::S�q��j���)l���-�5+ ��A�KP8y��-1{����;^e3F3����u��"�7>)Ǡ4��[�O��<��s)X	�셡 �����o&��$_�i^�g�}�dD�艎\�#��J����+��S�"@!�mk�T��Kx��ȿ4�"��5�v���z7��b�����b��֛��S��Z~U(�������$��d��x٪��jh�����~֌�D���-<�J�[,�lۄ�}%!7܅�M:�K}�l2G��V�R����+����]���=N��yz�`�z���wĻ���]�$��7g]$��[�O}���o7��-����P��  NXFЦrZ�D��7�p�#N{��<�sпL��o������O�wo��ۣd��W��ዘ�'���������Q���G�H���yƾ�%���d>:���.��`�78�n?:Ӡ';�,h��e�PU���;����5����j9`=L�̊_#(3Ԣ}!��5t�����N�h�xI�DqNTw �B4�M2/U1xh�7�$K�9�F��^�j�`����z�|)b9wH(Bq���g�|�.��Ś�	k~2��!a�lb#��U���.��_�a80#�!��ߟ^z�H��']��熗:�UFo-��	H6[�J?��H�(��}�ܲ��l�E�-��<"Xy��>,*>$�����pZ���,�L6�׾��s��j�(����va�S�o�$��۪�rνU� �)n��]{<��9����#vM��Ew�2��
Ƚ���#����L'�lb`:�<���=�(j~��r b�b�����jOsH�S��-���t�b��d¡x�Z����NVA�;�);XC�7�/~ck������=J{�E	�uKf~|�W���n�!Dӓ||:��L?�~�WoU���u�J��wPB!/�&)��[�t��v�H�����L���P��6��#�G��O��-7��lWU����oX�e�Ժ&,֞��|�)�|�6J�	l,�N���Q�o�;�F26���ب⒜�"*Mv�f��O��&����#6�=	�w�e1cB�4��Ij=�iM(8-��|�l�Y��׶�֚ιwk�׫��'�h���\���\⨡��syVi]��E�詻>�%nFM`%;%������{��7���:�y�*�Vm����گ�/�]�j�.x���܌��#AU/�@3S��<+V��!��~��-�[��u��3���SQ�_Q�� ��u �Y*��~������}\n�x)߲b]���U̓��Ia�Z�ZM�\��E� BtX� ���-�^���-9�IGQ*z�;s�E�ՀNmCZ@�*�tFh��y��r������m��8-=osv3�{C{Z|<��4=��<�~����N?��]�w k1��4�0̕�&��p/ǜ�5���p�(��I�mWqe 5X�
M��r]8��s�I���֘��۲x
�%��ؤo�P��1��G���Ά��
��XUN�d��;�(d���G޾���j�'$�jY�gď�	 �t��{LVk��0�rsU���+#-m���5�xdMct�@l`yQM�1w D-��:A�]$�v����O�!j��4��H�ׇ'
��������m�Y���������:%��=�O��[Z��d6N��O�J�|��T����U�������W/�ş5�ԗC���x�ΰP�����F��������G?e���&�K�q�~����+�.����dc���=��}�l�82�����>S�/hgn���8��h��١00üG�>��=^�y�G�����s��������]>BJj�H[l�� � 6�XO����?%��/9�2�}&v�5`%j;(��K�e�A˓p����b���
<"P�5�!��R\��o�/4P��F��e��@�(X��U-c{r'f_;�n/)cZ�q�t���n�/.�gi\$��ײՑ��kj��")�GI���4�'(,���r�G�M+����qY�$����b�yE�W#xY�ߌ= ��L�����k#�ϣ�3��{
�l��W��Z�Q��[�B�a������W�{��o���ߤʫ�共��˓x#ي-@%��T��K;EJ�3)wJ�T�*"F\\!��7g�����u�/���j%��"��ad�R�U&���-�^�>��βb��ħ�/f��B��BvO�fIO�
�6�WSs�+��ۙ`͡�I�A\P�STR�]i�����t��� 2}
q��"ho�,_�_7AP��Ե�HZ��3��R�e�yt@�q�D�e��N`շ=ԃ��*-4]��e1Acw4�#�
�/P�L��>!5�v=Ay���J_�ޏ��-|mX~v�	&�'L���ظNAI����n:6���T0�a�ܧ��0��f/ ���#,�Z�ݍ�mAB�>_�@�n��q��'�����'5:��[Y@/��[�48��-��D�=�$��nĆ�� ���9%�R�>]Us��=�WD��Rۅ޵P�sv �Aw3y�ke	ܩ�E%jQ��&� V��)���2�h)���*�g��G�� ;	��J'�ԑE���S�^���&������v:���3F�B�^�xF����B�W��{P]/f7VL�k���3DAŲ��ŢV�"�q�Y �~��c���$��dW����:v|Կ:�� ,$M�����:��O�xC�R[}��)<���#�ZT��rqRf�o��A����Yv�n�3A�7ʃ�H��&=�hh忳�RO�E{1:zSx)�2�1NB�2�JMިiA{���sxo�W��9�R�jX��s��%%��&rpU�ZLh%36�����ʂ�"w�WY,H0��F��/���`��y�XĺQ ��Y|#���ïb`�5�%�/W�v�Wt�m�*�nԅw���D����M�!r���nN̌S %���ݧ�;S�T n�8 5��x�k����'���[�.���{�{Hm�"S�YB��ʣ5٪�	�h(l�zDy&��Y�#D[0\_���6�n�M	e$��]Ҹ���(.s>%��A�v��i=��W2�ݹ^lZ�IҌ��F;%?����Tmo?�AW�����:+��+#�d�����4�4hw>�T%�7mM$��Y��Y�̰1rIg
��<=�y����bJ"Iw�g�6��f �Fc�[�`�q8��ǅ���kŋ����7�
E�ER�k���r�b��U�pk���('�H���=��/��<k�)ɫ06���Gv�$қ�G�`lc��Ԓ�t%^w,�
�N��f�B:����kt�R���w �{׋[�o��V�H��$"��)�7`�ÿ́6�B78���Ā62�ؙf�L��^��_�ǹd�n��p��B�s0����3�m+(,��hU�?�kP��d�[?3;C�z��kM���BB����b�ᦤHC�-�d��dIa�T��D�q�V�1�{m�'SY�{�2��=#�!�״ J��kg����w�&�%\ҧ���pS��&u�r�B⥱8f�5����(%Zg�`��؇�b)Ŏ�;>�u�&+H
`_�L�B�5� %S��tBϥ.C�W+ܻ������2��E�0h��*p��3�ZL�Q�+�@��H�R��H���v��͇��d�55$������b������_a��!ra�A@A!.��_���%�%X�}Y̽��@(  Dpp����g,X��;x9�	K�vhYi3X�vϮ��?�/5적|yZݬE?A!��^���$�M�Ŷwb@9t)��v �=�t���ް���� �� ~,uQQ�W�vԆ�<��.Yq.�~�)�N.���5[��ƬA�!-P����x��q&���1'���.��9;q��%�~z�z!��c~��l�Аa��M�A�����R�K�P�,U�y�	Ǉ�۱�S�I��z�9���7��uL�e�.,o��z��`�����z.J��_ϳ4P�Z@�8^�d8�LUn�]�k��	,���I��׵��-lǥ)]�-�*���L��U糅�~?���-���It�!�u�lz�:���a��]���Ģ��5X
K��&�^b�����;��}�[��)���F4�Vc��L��������r�e�8
��Cy.T!@���eK��;�����g���w�`L-d�|�]a�Ls�[�����<1ٗ�{�#�sj}����r�J�p<���8��uW�z�&X~�p�# �y�r���`>�%SVWK3��1Z���������K�wEo�P�{�8�S;��"�*ucL�x�����؞��l�|{�$L4O:����+�`	`ֿ�Ҹ���y~�IېL<T,�
�C+���l��ש~C�����IT�i:}�hάj��/a*�B+�g>Y��3���U�D�ӈ��U\gƔ֦7��*�|���X�߻��I�ڎ�y����l��\�yI��$V����������j��4���I!�g��ʔVpN|@�l�+�z�eH��?�n�d�\�~�N���3��d=�JO�lB�:3�"(t�B�
+�T��S�R���I�Bfʜ�����%�1U�+O�@����>Nēr��(]��L{��#,@3<�A��-�W�a%jM�0JE�U��f�	�Y���e^�>�R��Nh��������