��/  ��s��u�cx��/���E@>~���UҠ��.����y���7�I�Dy��Ȓ9���.7��r��
"E���T�rЬ�$�9�i��+w� m�l����9�F�T���4�z�ӥV)��-�7/��!�H
�ō+��fyQ��ӚP]��ud�m6[�1
�[c>�m	���39��V{ ^i���E�ቚ���l0th�*>�IjOd�ۻ� -�n�Ѳ	O�EM�%�b�v�W�P-Fe�MV0QS1�{�tP���e`/4���鿸��Rd���{ѩg�$�!��מ��8��8��*vv� �%��b/:�|��l����3Jf��a�"���rj.�I ��0�!i\��6��Xl�˝,^{�#�|D.e~#�P�J}�Qkx���>&߻$& mAs�~����q:�4�L����v�U�B��	�}��̈�|�rM�t�<���k�F�� Z�J���ʒq�W�ԒgFlH���l��q�Gb�����+�r&���[������M4Z�Om�IT��-K+�F
�&]�P4M�W�ʟ�u��jYw�盄N;_�8_"�#:�������mb�;�� ��J/�"�}�y�}��'�?�A�L~����Id�V�A;�9c�̵g�v瓤J��uV��ʳk��hN@9�V^�QHr��JQ4� έ���4>+�>��&���@�"��/Vq�㺊��9��0ܐn�C��s��yH�*`#G�l8^���+�>��4#<��=��Ʃj�,p����v�j��u?G�8X��sׁK�\f�7۶T>D%j��r艌���ฺ}'�Q���N���c�03Ai/���ͭ-�8�Q�u�Aw+Ռ��Y����.ż�e��u<t�pf�<��{܎V)_�m�G?�Z��Q��T�s琳�鲖���fH�
(����n2�@Z��Ϧgҿ_7�w�D��)̮p�B�lKB8D�To�;�}����cSW��ԚwӒ��{k(Y��G�J��|u�ܻ�c�abS��Xւ�%Q);��}׃F�סD���w8���"ک��=��_�i;��6�7���.X@������-��%x�v[���2�Քg,�k,�-ɟ��;��N��Z� ��1Li��d�D8�E�����;�!�1��z�Mz�V�_��A�#�3�|���]���F��ë_���Ln�Q�pn���fD����>p����Z���,,��]V�AZ��F�n'�����	�v!���'�<CɆi��r'��I�ι�`��:ܣVbE�(�q�A����7�����c��k���� ,�?�L����X>{�]*�r��L����fEh_��1Iﴋ��,�4�%u�zk��@k�[��yjW#�#����b/D�瓿@x�L�\����T<"�j��O�m���)��g�����(l���[�^����fP+�tH	^)��ncZ-�Vi��a4�%�x�to�)��h=�����H�x@��k�Cj�Ʉ�U��a	�
�?��HSo��x+M�TV+�T�7��υؚ��Ի&���g:��9��{+�M�.�����۰�7+U�����$������~��V���l�y~ȭn�m�V=X�<�"�rj(뷛G�iE퍳g!_8j#^]�2���Jf��B*tI����5��,��!m��}�Ӹ���2�1�MҧT�����n%�TI�.�-�_��Lv�/J- �Dg�G}Ƈ�K|�ΰ�+���):'1����\�!i�N�� Țp��9�9~��I����H�`vO;���rli��ͦ:_�;>|z�O�@[�,�f��_Č�R�u�񮒨�˨bD��|/!1u^᫻Ԙ�z���Vj�����)�o�'渪��ƶ�����s�7�L�,��H�������.��{Z����L���M��M �U�'Eu��P8
�`b��d�-�q�`�w�ĳ֪����pB�Fe7bH�������~�^��w� �x��,g�f���R�P�h)tr��.^�>|���k�T��+��7����9\�q��O�)Uyu��w޹O�@9o̷�hN}?YԌ���sݻa�:����{���������ݼ�ѣ�b�������mi�[���-8��ݺ�.�|"&�r�V�3.V�Fc%�P_%�i~.��.�!���S�Cꙉ~�N�yY5��{�Ј4aɻS�E�lx�3!���tq�)��}�
��¤��1>���t�kP��I�a�<��I*x|1\�1�4��9"#�����hJƣ�s�!e{����	��$J�[�v�v�����R�{����a\k���rh�������
4D�6@Z4���>��[������z�HBR��j�fL-�����6���&i�:>�y�pF�cvJ��nͲ̂|7"Adv�Vjw9���]���qf$<_�����=2��dr���������H9Z��5&B��NZN �&�+Vސ��̘�o.D��m������,S´���� l�l���4��Ӫ���a2�c�ݻ F��!n��Q��r|�<I٬��)1�i�*<������.����ü�8�kQK8��$k��k��ۧ�Ȭ��3���Rq�gS[�m͑3-e��K�+���u��̘�sl�����W��H�����Tn��=��(��D�Si��+�=����鿀�b;L����w�Ϳ�䓨��a�#��GL����n5\|�M<�y���t{�������IBu,�=F̮�h0)�o8�X�� ߛT��Z]��⦹����R�����=��F׸�ȹ6�'�x���(�n��������ρ����E/�������\~y~��C>�����L⤠�^եq3ҔD�ٶ]�GAE�篎trt��f�`�T��sK���?���	�{����q��Ai�j⎋���%�\�m�쳠K���@Y�Q=����3`uO��;ۥ�2�u��7h� k�4C��f�UJp!�;u<�^٪����Jn��4��;�� U�9�أ���)�.�/�㣙��D�A�+q�v��7�ې7�3憑@j���xݲX�����q�f������`2B�����!�~S�k�/2yW3�>&Ui��_
 �5���V:=�xi�DP��\�B�����ZM��]h�]�k8N ��ԐH���ܓ�J��8͗��D������nj7��͡D�e�����(ji|P�Y;�ij��[����7KtH�z��jÁ2�ZoYh�a��O7}����W�Z����M����®^#�V4�E`-��}�"�76?]S�m���.��RV�ˠ{Ks{�X�q��O�t�@6s �:`⠁�aY�����
X��F_�:*��*sZtM��� �_�be�K��	��5�o+o���:�83�����|0�;Uܥ�m��]����m�8�O�á*qN���?\�����F���Q8<OU0��F�`��?+{l����S���6G��>���;4~0@;�����&.3yvKB'���p��V�K�����l���A*d#��U�[�z@G��V��٭ �b�����ϧ��-"��sbv�l�t��/N6��%Y�lWbȺ�e`}yI��{���v����}7
u��{�Q����1���1�^x���\W��r"(s(�� ˘����#xI}���ߕ�׭��b�ۅ��a^�Ѐ8���mkz��;�tY����B��$�\���k���(��ɮAE�����IM�[�x<��[�:iޏ��O��d��q��U{�c0�a�	J`�nMM���4H����o��ey=`./�M��l�9otk��(_5U*�hK��*X���Y����Z������0ĝ���D�@!���ad��,/~@u�)�qܥX���^�nd��3` Y9�݇�ݔ�I@�4��B�13��+!C®��ĩyeG�~����V�p��cφ��(#��Ď�I�SI�]�$�O`Ne�'>�!@�=�����9vj�h7F���$���'���>��U�SED�F���1:ڪ\/�~��.]�k%B~9a��?�����
��/�x��tM���M��vYOA�Ԋ��$<�*L-.��0�c�^�m�8lB~n���K_}�<�3��(��������$�G����"��"mN���n�Ie�gr��i)�,&Cw�{%�� 6\>�(�L�,ՍX?�p����Z<�+�:m ��N�!D���v¯�=eD�]t3�]M6jH!��.�bあ�t�ʽ\�Aп�m<#Pd�:�k`��*�Y�ԯ�~��S�0U���������*͗�6�	����5�2��vm�8J��e�!#��7�y�fˀNf�t�F����(��S�^�~�^��s(�s���k��b,��V5�/��4#��j��Ʒ��P��n�T�{��S�B	u��>l�l��JW��L�ۆ0~���r��ZA{�i6}��g��`�����$n,���C��%���(�J�Q�̎�ŷ�/?��g�^2'̹�)ƻ�2;���<u�����-��=ڥQI�A9+���
��p�*���C(��	ɦ�>mO�k�v���F��j#�Ƅ]mQ �>@G�e����D	����^���#����	���@<�<��z뭓zH��D~�äD8b���|7��t�h�vHv���;<���5?��f�e�|�wg���gMD �����2�լ@�P-�6N�V#�l|�\@r��-�Ћe����`�
�gu�'�AVR\�%غk1Z�IKÝ�?�u[8E�{=�%r|���4[��`+zb���#�|gBS���}�2z=�@�<t��%q���r�Z�u�
n�������tG�.v~�)լN��|�-�5�LA�(k{%)Ep���x���>'�������EѪV	�������c!�a�+�S`L?dGʵ����pq�N��;O��'|���z�ݒ����0��ӟ��Lu
i�1�DCD���_w��ҔRowLyW�Nl-�s)�T|6����B�$�[�D����0�mE�e��5��8K�D����;Y�s�>/��6�o1���Źk)L�4`�Fȶ�:�e|r���7��:�ϑ�u�P駺�vg)u�[�1I|]�{�k�0D\���?V}���Lv
��\ޛ�n���~�H^�JD�;��|iD1�1�K]e��?3���İX��`7�vI��}br�H���H��-R�|NWϖ�Cʶ��7Z� -n�{\�x+��.�#B��'ſ�me��S(�h��
	_���XLg���>���ǭ.����F�/+�Y�՜_�}q�u�LT^ˇ���xZFP�C�i,X��z�E'� ���M@?.�8�aYZ醀5m�w�����8�M�r��yx��_��-K��D�~@n�!�_w��t�@�6[�\'tF5�WJ��v"A��Re	ҩ�{�7�uۚ���·L!��ꬻ�z;e�c���,���x��� ����'{^ ];Q�׌_D��4�}`� *ٞ���j�k}�V�z16�T\h)P
�р]��+���3|��/�ŗ�e�4��4k�f%�5	5�E����J��+Ӂ�T~�f��k�|^��_��$�A��u)���LA�l�-.#O;>^��̋���0b'��:�� ���WABtc�9���
}�qc��{Q�q��{!��6a�
�B��[85�L�u�wz���L\�P���8�-���Lw��l����桧n��Ǳiߛ!��@n�>��ih��g`
���9���;K�����e��IWl�'ĮB,�݄�ЙR�Hް�Yi�I�>4�=_7���MT/�ˌP����"6�'|lx�m��Z��� 1��]��X�Nm֯ (	u0}rf�{8Ł��q��P(s�������k��Ah�@����,�ak<du��=m��Z5P��M$VnS?���
f����Ο-i���.�n�i<[b$�Zʙ�8��B9��|o�(�y����RɨD'ۻ�	~O��_��t=M��}�Cs��@c/-7�Җ�!-�.!p&Ԝ��u��X��3��?��1� �=��,�j!�@��.���y�+�qő�w�8��O]V����ȥ�ϵĦH��9�b�,�wY͠&a��@�b��n��ʽp���P�n;�'�� ES,��K���%�n#�	��[�u�U�NP�2�4�7`��r�u��j�:�#��>D/\$�ǿ6�vE_$�6�~\ln ��4[aK�0�$�r��#~���Ĕ��G�Co�t�l���d8���n�I60��v2���{�����pΰ=Ԩ�D�d�s��_�
����	�WW�-7#�0Ë�zL�O^U����O��ry�]�>�s��- n(��RxP 8]^�1�K}n�Z��+bd��P����֝lT1��)�����F�ʭcmV�FjT�l��u�j��#m�����yPJ��vYQ���E3NC���	�����C�W����tU!0gB4_��.�º
K�^J9|3
�Ѓ�ѐ�4�%29O8���Ѳ�X�z3���^�Z�a͟/p��M>�ꦑ����bSf�_Ó�1Mt�y�w�е�1Z�n5"�܉�g�_�1'�<]m��%f����'=�=�Y���rq�τh9���������?�R�w��.�r���ub��4�N�&P�Ed�,��j��<��)dI~��8�k�g���槩��$��#��a�����?����y&��e���H�����������P�e?<��&݀ �Ks�B5in�J�M�t�}��3���!�f�s�߿!���#,k���9�\=Z�]��
�Q�r��:���fՁ�d<�Ź6L�zʵ�Ky���e�<��F�mr%�w�;-���Š%#n.z��n�P��#ږ���YA�����;�V����.�;%k��.�������^�̈�������Ue(��{x���Y�-$ƚB�֎��Ԙ�h�efn�2�N�f�����~Uy���ɀV�� 6{���Mt5�*��{�2ou�\y�����v�4�P�[�.M���o�h;�R�p�=K��<�&gpF��j�UX��ؚ�m�f���㱁�T�-<a�EMț3&0��Ӿ�r=:���J?ꥂ��Fn�tGB�.km�G�+zj�5}�w��V/�;��2!�o["�M5^>��H��n�%�X���L�;l59a�u��,#f7�����?���3���̤ 89L��v-bI��!5�P��`4�3��_�_�w���F'���N�~C^�Y�M����	�t�����ւ��1!.q�^Y ٞ�>�����O�Z��!��K�-�~J	���a�='6������J���$�(�n������D��"�c�;�%xi[.*�<���+�:�VEE�A�Vf�t���f���>�Z�,��=M��^I	'|w����6�w��\��k�v1�8��n�+�UR�<?cV^�sN$���M���4���b�`<��ϕ��U"��k��X��WR��ؿ�S��K5�xfE��3��E�j
�<��Ƣbش��W���x�B7���>���<c��|w�!���9}ӄLIo!U�Y�����xn��iF��Gf�H��|c|��-�U��;P iѫ2I8�����8�T��G�5+bm%.�������R��P��%�oCk��ld�'�dDGh��J��� Xb����M?���]�nk 
&�'.>\���k��6����VYhn�jǟ?̼��m��vN̯>�$&堹���A�B$ X��"����\Ű��� �G��mJ�Vv�omqG�J�54�KN�J(���aY�n�&4��l0�=C`!O���;E���z