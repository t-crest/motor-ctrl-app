��/  �W�
m��x�d���sh��6�m�9XN���Q>�\v��������))��O�:�]����B�Fү�����)������YURCw�Ѓ5|sf����WF����1�c�М�72Nl� ���YA�g+$D�ݏC�F���Z����,�z2�,�^�B�Ra��?rz�Ҝ���n4��Us$IBE.dL�0>��Ѐ@�\
��:ppզ{ 6o�br��Ҷu�:���9��Ԁ,��r��'}����ʢϓ+�,�u	��If�SZ[aW�M�W��������blT#�Ѻ������J�z
�R��d/8X*rT]-���`�c'f����d�;����{��~4�i7����|r�����~��i?o�����֕W����q����ܺ^�*C�k�hR��H'�P����g�-+w-�Vvn�E�T�6ӼL�|~��{5.��p�V�����b�&����Yw�0?�LC�1Zpڷ	(p�eVPL�[��j(P���}n۵�3D�s�_
�"�r�ؼg4����Ua�uN����Fʕuͫ܊�}�����t�u|��*��v�Y��NI�ը�ݴu�={?�,fو(��\l�*�Mh�5�������^�:�G_�N���y#(ƚ�>��ۼ���s@��z\�e�V���Qf4�ԅ-7�;r����9�A*�m��mW�e��+��F��<������Y���`��j*e����|%�J��b�g��	��{�c�E��Nԙ~�Y5gL;�ac�?u�m�̠潄�m/�Z�UW���]������.4������޽RL���xa���\����(b�׉���U>��W����%	������pE��Ŧ��*W��z��m�Fh���Bm�~w7�P��{��E���ꄵ9��%�&���d�v�6����FH���$�v���4<�,��\���U| ps����YR�z�
&	�����JD�{�S;@� ��o��O�M�j�wp����!��n�Ij@���F+���|bcO�@����q�EdO%n�{c��C|�����+N �r-���??�s��V�MB��e�	�ŝ�9dO��5ӗ������tJ�YI��\
C��F[[��M��-�`���Њ�_�f��2J����u�����M��&_�^�1";�K�\���z_j�����#p�ƞ��p�X̛Bɇ��9����#��JE]R��Jϱ��Fo�5+�4�.�*�]�-��[�a+�P��7��;�}�m�S��GH'��B����=�v����)A,������ز�ǡ������N٦���c:QD���f7�nF���NDKɉ���+bQӛ~��(������q�]�>�+ϊ�OP�K��/'�]U(�/�|�p��3��IC�^�0f�fz%9����,ZTS���;����V
>��2߸P>bpu���[��=�doI���Kǲ.��ʳ��'��m	�·��z{g̋��\��4s�x���/�5d%|��+rT�d2�;�)�ͼp��M������H1���+���E�x������UyL��d8���m�s�����X+97zD�Q2鱪p��Ķ{:a���!>�w�M��ָ�lI���׮��|�'e�L�+�y�����+rE��~���c��o\Bc
:��(��sy^?�ȍ0���`q��	��F9񀚙�H'�< d�H�_˽?�Φ����
��G�Y��j��D(�b�ۭjX3
H_h���*
��o�)�C^�Z��6�ǂ�a��g�g%���{ۇ��:�7�¿:Ho9�k���uc���j�0��^=\(S�?:�5�4�,��D��-K8�ǮS��g\s��ΐ9[�(R"a�y�����c�7�4'�t�p�`�d֖�"���j���(���_QTMbxĄ~NDd����#���Ϻ���\Rf|S{Q��[��T���8ۦ�l��Z�<F���,�س�Gm���hx����ԣ+�ҝ�L�Q���S��mF��,4�@�*^Va���7y��[̞���ѿ�^��"�`6�����=X�mV�R����!�l�}��~3k<�^�B�v�nR��5t�ө(��F!̟� ��)�kU|�!�Y���.�@v�,.W����u��K�s�C�Ӹ���G%(�Q#Α�D`uo+-���&����(�d���IզsGs�� S�n*��8�eH��v���06i qr��-���J�jG��|�;ژ�F/-�N_���K��}�XF���;��	�3��<��50+����f�}A ���%�G��m�_NX� �������N�����9�uF�a����IV���m��~���]E%�,.$�{zp?�_������"Q� d�����-좓�א3��
��2��h6��#���^fr�S��7ٽ/ y��#[������Z�.���77�����y���9Vg�"u1���Z����E-��Wȭ��<�p��D
d���gⴙH�����	-[+"�|�0���k��G�p��Jh���/���L2TQ ]kr| �����%.�hY����\UÊ����xu��k����XԒ!��ל�"N����$NŸXDsѥ�6 }_u�>��RI��(�ա�2�<����Y�+���u�����.�L?{��;�����K~c,�b�vm㙖[^�6f�����q���墣�y�\���9�iÂ��Si�E�*��t�	������ڋs�*Ox6�E��&�h�#L�Tr��=[��c�5�yY��R���������}^�X�^�@��
<���j{��4����Y�F�~�}W�c�x�X&���S��C�D��r�td)��?�夸���Ce���'�sz���zw%5�����w��+j�ȵ�甊p�XPn�'���Ŏ(l�?t�ب�)`4=�t���U��!�ۿW����]��wI�>���.��g�ڹ:n�HH��A�$�}���t����� �E���	��Zmʻ�j��G F�?<ߝF�-�D'��s�rR���|��ߣ�%�ob��I,STo�u��dS&9�F���ԚS��Zµ;��O�ė���i�3[��R�Ene��� �s� �Qf��}1�A=�����JĄ�߁܄�)� �U�D�}��F��-}�m�]X1��7!b��>U�_�4#��s����j�����W��p��(��Tu�9��|�$j>�*��} b�����n�x.˲����ڐ/�v�� �ƆL���$ �R�0����H0{Z(s=hc,a���W�P�Y�'��B� ������] �
����s�HT��c�cQ~R�m&�sȹ�9��D�����r�����j��v�)d59��ذ։0�\A�3�^hKG{wþDy����z��u���Z����'���/�4��#	��9]�ʛ�q*n�ſ�-� \���t��.�i���]P/�aI�N�R�d��m"QD�/����G� �S�0G�C� �j��v�V����;�2���hV@~6x��B_����Ūu%\B9��uy�8���C�j����\I�K3�*��������KFU�>�A���P#� �8��gTi����^ަ�s~:0����6%�]��}��˾x`'j�:�>��w������'�궽��;� fw��G�a`{$\�~A#2�`n���6Wx+Tx���1zDf�J�k�!v�2e�\��C�i�p�6YN�b��y��n��\�k9P�k{�r�����ݙ��(zgw����1����߳4
-�K�/u�H��g~����� lc�8��j���n�vLYZK��0q�S-�,���X�ԏ����������o�ep���K�ն����_h���=!�^+��7!aS��� S=�5�������ɝ�X��3}o�)�*�f
PÃ�?����L5�h��P�G�7G�,yW6�؉�#FX�j���X)|��y�A���ىf� �"���?�ԶN��F�E�S ۟�f�ڣo)���K�r�4q�
d{���t�x��<頜l&��3���!=B�3�0&��rӈ�]�l�D�ֻ�� �3uj^#���v�q�C���;7�#U�XZ�����;��B9�cP�A0�eߖE��ٛ2�B3�	���~�B�Խ_�;��i���.��Ơ�<�5)���}-�Q�<�����������zuX��s��jk��,��#z�F�"��O�a:�"#)��J���Ģ���u�Nn�0A�d+��e�U_4BU1�b�SX��;��� �ȬG����(��')i� �b�eB(g��.b�-GJ|�<n'�y}�~��e�$ ����}IM�����g]���#7[Lx�Y&�ּ��5=<:�;�?��k ^�]&�%�1�ۉ�U�%�ҀA.R$Zw&!=���H�g�3��p�ڄ�f�`�?"BT���� �Z*�ls�9��KxD�n���*�+I�bY_��R?(i��)�-�[��ԑ`;+�=Osb�{�������<_�	�x��`r8V �en���#�� �N��R������� K��f�,Pۑ��7���CCL��� ��E^�����,������U�LB&ȍ�љC�d9*Y����1J_V����?�V]���b���4�Τ�o��<F��j�I������a�J��)ۦ����H2� ׏ ���Um�I�e�]�=��x�&�� �	��V)�B���i����x�4vXf���Ķ��� ��.�^���@�>�+��Kx��t���x�J�ep��jP��pFԀ^由OK"�n� a/����
��F7}3|\sx�6��\���nJ�"�5�����rD-HD�jU�7 2{>�]���'�l�����E~#�Ӹ��[�y�J䧜�;ªXر��Г5.�\A�-��|��;�C^�V�Ę��g�V���4,�!��+��ה��s�D�K	��$s��K�(��L>ȊqP3scg�;=I&V%��>9��·O|�͢m���;p�M��
��v��$�I+� 4m �EHR=��9-�ʖ�����7�L�aj2:�e��w�t����@y�T�o����c������|�XM�q^�=�9(���n@�K?����R��W/��O�@��&��L�#��S�qu��33��]/�I0Jt�<L;��W����&��&	�T�܄F�hn�8��s�*���47I9S�f�����{�ӥ����n �!8��ИlRI�1[�~�?�����5@�c(Y��}�N]��-	�ۃ<w��k�m�h�>B�"��X��bȊG����t�;��_U�i�g�rY0�$�N�1}#�)��%�z�~Y�x%(1��p�&��~.�ă��GML(������cB�-��<ڭf�;��C[��J����=����l5�����Gt��Fq���w.�y��4�o��BQKl	��U>��8���W���޷��W��'������6UKU+N�ܣ�,
��k���ݙ|�w���|�$\��A���4aU�;�����;�?�JGnʕ���+����P��fR�}�#���#_������е��C�"�"���ƾ�¬(�����5+��n5J��������?���ֳ0����D�'N$5X�7�e��~���1�\�Q�ܭ|�z�m}��������T_����r���ρ
��Ϫ��zOIS
6���;�6j��������UDrP? ߨ�� 7qs��2�tԩ�1�s��_��~=�<*�̴��Z�)��s�Z1�L�K_�l�"��H�J�	�3�{��}7m��"u.��/�C�Y]���?.��㗞<�Ϣ8���i�ݭ}�3����;Y�}XO|�Om��j3����<Q#Mw�|~�I�_���>���f��µ��ꯥ?q���Goid�-$$�I�ß�|���:u�5���N�{��V����"�/
߁�����y|G��F�I�FʋS822��,0^)�~i��ş��W��a��._ߏ�7���|C+�B��X���-8������]-[.[d�����\�]Ϣ�	��7v�؞ �hu��~)?�H,�]��huS�ɾ�ذ~¢3�:>��r������)T�[h�	�l���m�"��{��cć�_���y����_D�e�#<���[jӅ>��ٴ$c*�"teY�P�E58ɽ*�t�9�$���jn˝�e+ǹ�/����]�����pc�DN�L7.ډ%;m��Ԓ����V_��ߙ}�Y� �x���,�TMR�J,!Pm/H�A�@��$�)�ȩ1�g����i�;��a�u]
_�s��V��@��N�yR���,$�K��e��.���@��L�k�7����FL�s�``*Y��R}�_�1���}	���=�2Y0u;�Ohb P{���d��2M9p�K:��K�E���j�u�79a�(?�C���;{�G)� �i�cs���6��S��ฦ�A���[+�b�6M���7�}y�؋����TWw�%��.�-琎Eѡ-���l��ұwG�4J,B���5���莈�$���ř^$��3�4������	�5��;-L=�Xڌ��ˮV�qD7V	�S$��;���h����O�؂���t���U�""H�c��So#_xr�
-���M���ܬ֝!;8  Ç<UI�~�C ؅��21ad�l��7pf����S�U�6c_Lx4�V�^�S^�(fGn�B[��g��4C��H>����j�q��N3yAf8�$ν�d����G�߭Q��ZDkF���)��_�eH�ļ�F6����"��־�?�z�����#�ܤ�nN��k�Dn�V~���}Ҁ�6�����x��8of8� rz�=B�J��0a
W.�9
�[_��/vࢗ̠���rT�����
�~o�E�A�L��ײe��q��O�Զ�� ���ѯ،Rq��~�{Ny�=f�	NڅU`'@Y����j�X���z�:�`���i���gmќY�+����d��8SB˫�[:�&�)r���DG�Z���/�h��!���C:�6~�Y\EN�-W#:ǅ���5�p����$	p���P��&\Jق�}�෋���� $�i��ת*1�PM5�����y6~W`\gj\�������h�k	���	�D��e�:����OԳ/��r����k�L��^qc��S�AD��i�|��i�1�O��Ti�����t�`1iJBP5����U����b+aV�q?<�{サ�G���oʦ?�(&�-�L�2SM]��Z��@�&�恴1�w�P?KPyߞQɞ��S%�ǁiZ�?�U��Q��, ��,���Sg�%�u��� bm������"�k�'��p��@��/W&����CΫ�+�p��e��ߤ���S&l
u��A������C(B�g^�n9�߼'��k@��q�[��3��G0�z<��eXj�RX)ϝסu��TH�*�7��Bi��=��*�(^�-C��O��F���fp*# H�t��rD���N�m��m�f%Ow������"��Y)��?��C�n]x�O#X*҅�Z5k\�9]� s�E$��+�e6�&|oB��s#8�=59+]R�_d�c*�s^FN��6��9��{���f�H�7t ��`�;���'7��:�n���'ň�B��\�N���M���/��J=�Y�jԑ���+ :�ʤ-�zT�D�S�s~�\��&׏�`']_���i�?vt�`�d}k,��+ ŋuF��������>g�u��W���CKB�)���݉	F�_�7l7�y��C5'��x����d��T��Y�GB�\���h��\:MX�0P�)���G��d�k��>X�����ڇ�`�XKH`è�=�b!#h�_�.x��Lm25�"6���_�O;2n0aP�T��M�v[6d�.�s�FL��\�����8e�����F~�n��Q��� �Z`�j\���`����MT�{��4+h�J&��.)�
�'��8�>n�,�P��Qɪ:o�f:�x+�\1��ɥ0r5�fC�M��C��Ҁ�j��.��<��0��B,B�<��^��V$ɟ���{������݄���w��D�v����Se$�����W-L�5I!�tmZ�3~/3����*�����@�Z�4f7o���Hf�%i&��۠����Q�뀇�YD����#j�"i�}����
PA9��T���:V�4��-`6^�b����b��,8%��Ut�c��A� ٪�m�3(��r5U������b?mf���x��|��:�i3^����X[Ǩ[�A:=:���ﻩ�/>h�M��$��ʇND��훌k�0�#~�6�=Ug��|:29-G�D��6*�c{b�n������,�Yo�����0�8�],$i,#K���\�
?���#n�>�LZ7_8@��(s����������&��-���*��DC
�OCw��ȃ��J�k� A\�������:�B�33^:J��k��Y��m��R�^"�nnZ��	���؃ɓ�~���%b��A���+�e�h������褁Y]P�)zO�Q�#q���M�tj����e�V�6kVi�&�U�A	��bjq����R�Jr�Ay�J2/���,�E/��q��;���I���^�	wxN�>���*ykH���׮�L]T�y]/�1����Z��x���4�_�>H���JE��lE5��!�b�a�F��m��+����Q(L[�tM�<-bY����N7�Z�c$�/ ݷ����i��#L�.�L�?�,�Y$?�/���G�Nt𨮋�k4㜘z�K�=:X忽74j���{ 2k7��>N��K�s�p\L
t��6�h�f/�(�DoMR�		��p���O����|lTmTj��K�~�B�r�*{�]�أE�'̧9�����w��r���D*�'�]����ŇP^�\��I�tK;|4+�=�Uݑ��7�-Ɨ�HxzRY��R�������UJ�-2Q񊥳�~
X�FK)�l�p����%���'[�@����?�R���~����f��5�S��(�p�M�oD�L��Q2]��|:
��(�ib'�xn\Ż`�V�����ֿ�,vr�fV�%&�txXA���Nt����QZ�q��Cs�Qs!Kn���,��o����Ѡ���#39�	�CHܒ�{~U�+zK6[�8�I�1ߏ��=M�!I�ۣ���}M����˕�>�h����@ֹ��,C<��cT��WSU.%ޤ���}�Z�Ȝ;7���8���0�)�`v>L��#�zH�;�\g�,bΩ8kqG#k��m�|*�&6�R
0�i-��ԋ�i��uH^�24��v9�U�v�`�gG�
���I��-��?*�y�^d���.9����4݉W��z���{�}��|X�^�B�*�'�Q��h$��Z|#'S!�KS.��I�ݴ�";���q��W)�CW�y���k�����Q���r9Ԝ}��Or6+W���!�ɘ`\+H ���"zVF�;ꯀG϶jjhH� X�%�䖙F�o�w2�����4Tt뱃���m��n��M� ����r��j�H&i3X.�[ܭ~�� b,�yZ��d���|%�U(䧩��4NH�8v]��Kd�{��	}�����v���\�=2�~K*��[�*7���W,y��m�� v�>����y��y	�>���g����g�+g�"�]Y4֡���R~8V�1} =Q���=W2��q�c���%�u����ѯ�|���m�!��o��{x����p�?��p�'�p�`r��D'-%��=���`_2��6󪫉����������[�`��y	]�i=_F��h!��V��ׯ?)*��/YKz?�k(|�G�9'f�WZ�T�$Hy�ɋLR���(�1�:��Ĕ�z�c
)"%\�� �S;�u(�Q�Q���[6֙�'N�sR"��J' ����O����\�*NԹ��˫�&��K+�E@E��L|m�a-TW��'�Yd�jY���	�b_�����-T��'H��dTeڒ�Ɍx ��Ė��R2�;�@�(�U~��O�f�y§0{���BldW��fį>l�$��WQ�\)�G�)�y-~)��Fr��I��>�ņ_���),WI�}x��V�?�����ɄP�-��~�����������Sk2,�je-��6,feڗeXa*�����Ϙ�g,�5԰�=+2q���S0��!�с��4��M�å�h�8�q�
x��v,[��@�%��R�ֹ(/�������&��dsy��g�zlU{$���Fε���1��^��ݛ���U�_|��
K���"��(�,X�yr�q�a�3�/�=~����-"y��jE ��''Æ^Ϸ�FHS{�2ϔ�u�ɦ��y�x�P5o�^�$�~�6�C��� �~޵�Q�g�lgW��.��|c���n��?W%MO�rj�Ͳmވ.��c����o��>Ԋ-��x"z�Φ@E�DYD{@*��������Ek��5�Gj��E^�ر�}��0��9e�k�o{�
���F ���3�g0ǰm�]�B���%�;���7<�G��T�`�q��<&u�t�wtA � 鞭TEZ�� �$(s���)�������s��� �,"�4��+7<v���6$@�dr5����w��V[;=l��99
%����ο�'y�U�9D�u��m�0�vh�P�W�U(���)jo	�'n�𴎉�i\�����.0�&�5^�z[�W���� �(�Y��d1�R���0RK�z7�EH\P5;��)ڷ�<��1s�m�8�Gi��ӵ�Ԡ��G�pm�C�$:A���1X*�@x�NA.莺*�9ہ�\���!l��a86#	K�ܷ���"C�I�T��v�с�����Z��ꊀ�OndP���.WVo��FZ�*�f��`��	6�5F�T���묙�-KZ���?�	��D���P��e�;�WR  4Wo����h9��	�P�2�Nx�C���=��_1&��'�m��c�DS����N���	F0��*iUesA��6x.P����j��}���ꄷT��	�L	/p�~�	���c�~�t��c�.{�A�!W{���E��XJ]��h�(�	F���1���U
h@`�â�����oSB�D�!���Y����;�K��Fz�%;�:�/k�Y��Cʿ��;�뜀Κ�tA|��� I�s��<�\׺�G�|$�$�Bc�{�_���e7"p����^z����3�������\�bG�h%x3O&�_6*�[0*d��#���k.�Eћ!�f�4$�s�zʉ�_�f�֞'��:e�����e\!�(>C<��li��F�}�p��Q��
��"R~7�z�������̬L�':���P>��iSʵص��H�x�Uݲ�P�KV��܇%��3N���`#��/��8����8㤑+�7�� #�j�0M�9՞-�/E�4��V��$h�݅�u�+_���'桛v�ѥ���<���n��KzYv9r�O�wЌb�'K���2�=�ґ}��)�����e��^o�S���
���
�:
�=Nݐ�Ykx��y���wg+R8w46�hf��J�G��οK��%^�P}���f��=T��Cƞ�����?9��͠�J~��ƺ_�uX5[��<�>{ڈ�Y�%�� 1!���O7&l��55n�Ap����(���K�L��\�a�Ш�>5��`c��p��ҿ8�%�
�����S���j�F��Q"�G_�F�G=��7�qV��*
�� ��� �D��H)8�:�$g)\gW����5�uW3��4� V.T?��X��S�����ZԠ�Qp�Տ�x W�0%��{-S����i���؏`Yn��԰��A��.Ŷ�P4@R�o�~5Oʋ��9T�^���F^�ׇ����WFA"i� ���5p><3����퀉��7����9� ��N �����F�L_<,c��q:$B�Ҙ�z����᥌UN��I<�=�ֵc�	�%���B���PL��J�F��eKSR2����m��D�8D����v�U�� I)���J��!Li�c
��'~ct}�� �.���0!~DꢄM��8s��&S:��8(6�՟O(��zBR}�%�8�-�M
����l�&�#�/�KZ� �w����"Z?�[�Ce}bm���$��׍����{�0J�O��� v>)��sS�����rj����3`�_
b�P�
�3�/w���(OY�3*�M'+w_���!�$�Z��_�� �SE�!�?���}V�j�s�Z1�S΄��F��N{;��w��(���Q����x�԰aB��R����7v-#��}�3F(|P-��N��П�ø�`���Bs� 1��>�ʱ?�/�۽'�S��0	�;rw�	���@�uWuz�x	����i�
6?�\X�2?����˟:�-�̱��C�é�N U=U+#y�A��]���i`�����2F�WE���G��c����'�^z�� 
�!�n��� %�'̼m����}�}���u��B�B����'����;4�t܀�]"-߮�*W�/=��)j�u��Y��>/$�Hj���eˆ7��9w~S ���5\16T���֑_�DN��
y��`M�2D�Ma�M��a��i"g%T�W��%�V�~m��G��g{���x6��zC�1���Z�k
;�<e;��%�c_�'$���5�`ֹ`S�V�1Mʹ)d�~��s��eSz2��;�)A|���z���3jX#�]