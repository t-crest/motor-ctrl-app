��/  S��3VQ(�x�G.���<AZ����O�Cm�	)�@�Z�*�s �����h�_�`�q�{��ȶ$T�}���o}\��3�Z��r<�ܛ������Iyz񄱘����&��+G^m'+"^�����)��R&P�$g���rU��d�DOiaٚ^��<�J	9�yI۴�:Sހ?�!��mbH3.��^;�b1�A��Y��7x����i~?��@�����Ǵ
�����^�d��%ÛֆI�.�����ouY�ʈoa����*,};�HT'V��t,��;�
$[���Jw�L�f_�߸�!�X���RRp�ڬ����+��2�͌���gǚ����*`z�����e���<��B�x��D�^͎2��o���� �4���a���f.�I:�U{�^���[�eߥ�@��V;R�p���|Di���3p���"k��NF���@ x�~#��T����+��5�/%�jl3i4���9Ec���H`�e0���umG)��S;@�-���nyL�_�������/n<^�#�TP��i4Q�e_PEϡ"��$V��#��K �?>�t�(��hO�+�/�I�.>y�)B}A�<yN�@��J�,֨���=�B"����@ )��{%��b���H�KAG���rIJX :�������ϥsa�B�e/^�ٳ$릻�����b6���&ܿ;}�:<ђH��jbx��+g2R�o�I�hn��:Vi�1Qӑ���[�g�ɳ[ϖ�����6��$`P�	{kJ<�N�H���q���� ���)O��g.eR�æ���MC�Ҽ��rɨ>�)N������Yd8LL��(l/%����2�<f��wu�E[r2!����P\@�s���ڿ��W�-��h�.w�X
�P�B�u�f7���C:��^�~�X�&~ŎfK+�M��;!�b)��q�$�S�Rd���L�k�o��h�'/���e>p�Hh@�#���{��Z�H�("8e��=�; �WH����O=6�^,���\	Ś���7��t��G�����6�s�s�ci�]�/ˡ�N��߮0��)��fz�~�����*�Iڕ��t<
j!>�1��MȪt���$�5utj���~�gN��"5��p�>5�Y��CC�Ŋ�P�ol@9Lz�Oְ_�J�3�،����6�5g�=y�˿�i(-ީ�u�t�2��"��0ԙ�,h`�A+�1���s��#��f	9Ԗ���D4�S���)0��e|m=_�,&�����H�[8�����-� ������f?�pR�lT��0
�:ynJH۱��+�*��h��z/���g�vM���}@�v��#���xl���M$�wIc�c(űp��p�sC�G��~B�M����ߢ�:�?�77t�]���x����t��o�������WA14
OZ!O�k&��nn����K��)l��)��)�V����<;qDz���KLh���b	�^v����@ ��*;����-���	s��;R�Mc_��1�ܫ�S��;���!�L��LTo?\`lG{|����I"�rK�1�����Ϳ1��� �#N��m�6���+�x�ԝ��\`�<}X�Ќ:`aC<Vb}F�Xrò5���e:d����M'�bۙ�VQ�L���'b`�����J���6C[a�0�4O/M�Y�PB���6�B%�>Lԑ��`��F9@k4��S���r�n�q��nb@�Aܛx��� X�q�����V��@��0ε�A�[���-@b%)c��Si~�Х���?Vp�j Y:����Ňz�����d}Vr%]IP��d
��h�|h�h�|Oq�##KH��2���(�I�w���I�f�{�]ڬ���-�{c�e�w���jQT0�Q��WSNу���6L7��Z��+)i	���>
Ӻ��F�%�AR?� �?�-7�s�(lV��}�d.��W���+�i��@�$��>�w�45�\)�Ys_�����Cаi�Ms��C%6���*����G�Ux}��.��/I�h�e*:�}n3'9Ek��;��K��z�G�`�Xݸ>�E�&�<��i�y�]�)�9����|��7V܏�j_�;���ò �x���D�yx/�dj3�u��YH�g���*��G�&�.K�K����#�����]�r�0.=�����Q��ӈf.�Ҁ����:���3�:�˅�����ч��#z��Q��f��fA��G���5�Wk�m�^S8�빛(pW�����JN~CBL[�s�g�Z�&�����$&��VyӴԫ,Vk�{��E��.���`u51��.�l�&�&�S�<%�i��K$���T��l3�D���|w��Q���<�*�
�E��V��)Q�a��Sh�w
n"J�BH��'��8~���:�)��"0E̞D��q���[y���S/}����ď��ӝը�d] n��H���"Zl�׏����.(ŤË삼�iEH����o$RH�ӹ��4?��ez'.�SR}b�Qؘ��o8��X�"�}�D��9a��ԁ9�c�:���n(�=g�;i���wC��$>�����ď�˵Q���T�q�'��4�R��W��k+[[|��r!�x/��0!��gڶ�>�IO;��f��C�H|�Md�"�%�]b�\��R\q�M�W�<G���v�_�^m"��~j�3���ۦ��8o���\w�*�-�ΩA �DStp���ՌY�9�ӏ��D@�ɟ�����.��'�[L!�F�����ʖSX��i�J�X�8���p@K��+Uf�s^�"ʒ^|U�8�)Y���)0�l�lS�+�&$�v���S�W�e������$�U�.a���r��d�8\��y���q	�!	v>Μb	��;��'^��2pZ�}羅#����d�n�f"���@p������	CڂbTt'���Ts4��טi`�H�͛��u�H��;��4�Y��h�=�C�B��0����PX>&'t-�u{��Z<�����-�'�V@�99~������ȋ�|�����b�V�����T�	�s�փ��øRVb¬*t��1�+�u�ggv�D��m�y���Pw�(1:�`�n�2uo��6��O�a��MV�)v�Ii�1�[,eڐ=�c �rC���&�+��W�H6f�j�r�,C��<.ɼ�c#���g-��e?$������>�e]��Eޱ�Ll��N�^��zF��t99f^ar��y����F��,�������I�j�~�񶂱jCvm)@�1Vj�V��p��DM�(.>.��gk<��3�_�/�e�,�Y�]0G6�կ�wq��[�� ���t>�̶���g�ݴާ����襆xB���Î=��T��s��(�u�J��
���\�и������r����r,(��qz|e�G�{�Hu���7$�C�sHxxb� 6�m�v}9H��Y���e�W/����'A�b	�o[Z� c}	B�}���H[P��2Q�j�=��W��#dRRN�:{$�:j@���7*<դԡ>�K��}���2�1Ӎ<l)M����C`I�%�~b��N��fK�W�J���nP�i����8���% ���}26�$}z]�M#���᡾�F�fM@��o��S�"5_�BK�lr�����[�[W6�		'�l,�3�8���7]�&}Ĳ�]�����f���4݈b������ 辭p����D�����klW��4��m�-{��j����]M��䡆4ڬѷ<2lm�k����e`ԙ�/���	%��7�ϼ�0��x���W��`.W��q�5���D�V��jg���Fo�U:���s�x��'�u�=.hv!�ӝ5)�b�{�h?����\�J�a��?��0�ԋŧ�:M>��Z8���3�I�L35܊%���Gų�R�F��8�Ṅ���x�R��Rd.A��K� h����0	y�,#�q��>���_Ty����U�P��Ά<`@�~�At��:]eB���c[��K�;�,�:�d1J��GX����i�k�s:~5�x���r5�+9,6h�L�C��d�O��w��54Y�6=�1Lm?�x�8��b��+s,�扷h �p��gv�c��6��?v�Y��J�����1�4��7v�uH:`�V��Aj*_b����6L�`�4]˸>KO��T6�(<����,�J���p�*B@�W��Q��))�R�?��@m���+|,/=)�L<��X������J���w����`
�-rD��<j6�
	�fz1��Q��ߟC�;'c3�7}����(��Ԓ�pa�8n>�F�t|W	ʤ*�|����^������\�b$H:�ີ"n�a]r��t	�j��)Ϥ\�p�l�q����n�$�������<��'Bh�<Cg?�Jy kqe���`)��L����-�ⴇ���h��S�Ib�<y����p�-�
9�cm�K7�����Ir���+G*?B��vL3��p\`�O���N��t���i�7)�j�:dW[���RZ��9�fKZ�,F=M�&]+�G�oγ?i�U�["�%�Q~��fsz���Z�������Ìf���np�*��~�E�i,���#�Z��;�R�k�':`�H���biU &��Eo ���<3m�<6a�c�#|�/
0�w����A=	�m�wT�O�Z�2a�����
, ���u���sB�ΝO{�v�/*˒_��)�a}j�m�����z���z�]�Ť{��AKF�~�5���C��%*}V�D9Н�z��,�����[��S�I��NQ�\����rـ��gBK����}��Y$5��c3�r�a>` �=o��:�@�"'�v؍��I�N3MKWi�2���>�r���{e��[�\�$bK|��Z�3G)�Q?&y�+l	�z��37��0H/ԤWʭ�VN0;�}�*$����E�g=%��D3����W�	��E�C߼����£1����j:�и�0���T�2��X>W��p��6��0���S?R.��Fv�-����(�ԺK�1MҮ5��b�; �D;�O	�E�Ni�2L�tC2��.��vmY�_|�fY��7���c:>q��ފ�LK4��U}%z�L�K6ϖ��gK��Z�4�کkK�����˟��H������[<,%&���~�:�ӚŽtB|Y�>9 쨉�_wS�l�)f�T8�u��I�úC~�ǃLB+��WsF��y�s���x���3H�y�\5���?B�I�� 5@� S�T�>f_P��g�Z��	��`+��*D6���,gu>��vbHk���1IBU7I�{�~��#�j����>$�jZ���{�҂�H�>��լ:����������	����9<���otD�����yC��I�#�d�N���q�9.��D�u����2���Q߬7�8�Nk�K�@2��4v�Q����X�� ���4��S�t��@�L !�隣iQ67+�o�ƚ8�g�3�:�E�_;���4­���t����ۄw�;�Dj��Vnn7�$���a�,g�+�Ȓ0&�A�2�,�WE���T�\�,��)�:�0ku��͈�J^���X鋢��=�:;����^��C(�۠��,$����R�z�9>P�N��� ��t"��
C�J���s�#Du����RMum��d¯�L�����'� K��``���c��5�|5���7�|:[0����RǤ��FN,�8z!���T�O2Pװ^P����u��6��1��0�t��(hr�"+�+0�����>��Bi�����-���AYi0�Ip%Y`�����kh,\����H���W�	u�����i���ʦ���Ƥ��]|^(G�y�F�3�0��!��u|wpp��©��!��0=��l�H�?��~��%�� �m�8���odJ���Wh�����'e��F�O�'RX7�o�jz�6�V��q�9U�����&�(1�w�����f�~�m�KZ�=��>�(�{E�0\� �_�j5�"�{ç:�R6�A�2)����f_G�;�}K�8 )�1=6@YyKp{ ��g�ؑ��:�:q����C
��8�ԋԠ��ԭ�B�ͧ�K�!�)S�R�'��@���쯭����M�
�>;�)Y��F,���$ʳJ�7�ބ��.���9�k0/����O�{?�'ۇ�ޛ!���	�����l~y1�ͷr�d��B�C��"P���`O��"�$��ۍ�� �AX9E;Í{��3���]:.�����Ƣ�w�h������RxA:��Z�y~iI_�F:���E�'������G3�������R����I5p%I������d��=BU4v��*&c�аL��D��prm�U�iP�n7�������8K[oS~�+񧓂w宍IQsua83a��)֌��c�����Q���)��@Rd���^{�x�M8m<�e�����bC1>)�w�Є�ˠ��g��j��v�ئP6::�Ra!������_���01�b��%nc�i���}���a�SfW�d~+�sI�b�HWGj/`k���ƚ��i.���Q�HfJ/�y���p��bl�;;����u`{Mz�R��92*���Z1n�'�Rj�����, �p��i��7t�5�菢1���@(�ϛ(�b�Ǒ�q����_�eP}�sRC�)�9R�O-�6��g��?m����y$/��su��Tv�٢��4����M?�p�$��ݴ.e���J ��1�ړ�����U}�y,���-lKwmi���j}�٘8n�?m���H���"��g�&�K�08/�.��x�Մ�T�b ����;a�o��j!��LXȒۭ]ϫ��*���̳�c<G�A,oG�y�%<O�s��f��z&3,i�ѿB[[�Yø��R�%@�U��x�4���R�	�?/n�-}��H�>@�x`��w1��>bC�C��+�:G=�s�"%�?=�R��DP6�ϊZԸ3�)�$���A�fawy|֚�?����ۮ-����v�	 ��9]t�`A��I�	�Q�<baniyaT�p�ZIlg4��F�zP�$qf�f�:��6���ָD��f�F$�Vc�seB��k���¦擯�(� �*b�ʋB��2���Ž�������d$5}�)�q�3	L�	�.o�Dė��dL��v<�:=������B_��E,Q�l|�5��X��%���;RQ�6�I�	A��ܭ�H��`K�$�ֽ%i��*�P��k�"PC2�8�P��/��BUd��{��c}CD0��I7(�M�a�0lYm�!
`�����әi��[�0n�}	�[�e,�*�5Ih��Wڪ��,��E��Mtѝc�����N�*@��x/�z�P�q��HX�ln�ѫ��N뾶�������������S��	�M��y9�{H9�xN�y��* � ��!�[=�T4h˂�ZF�آ�e$@R0�yb龎>ڲ�f�v�:aV�vמ==Z�E��B��E��#le���Ӫ:���C�p7�WT��I����~�at��{�y���w8�~�ܧ�oc��?,�.%�7��@[˭U&E5{f+�E�k��?r��9����Vh�5	���0i�ej���-G�p7�\k�9�7�R"���q�"�
W�3��v�r˪�4�J���*_U�[�^�HL�|�&J�h�8i���} ����zވ��+$��,�M�jf�F9�Iyܕ�ܻ�$�*5��'�	rs|B�K#:?��/��M��ۘPK��̎J����Y�@��`()e�qxK����x�;((�����96�k���g��f��4��]̥�㜒�I�0�b9�q?l�!:o��2�F�G�h;t]KQ>����S(�9uDD��9���i�����l��K�xL�'��x��E������x.a�@���X�Z2yq�z{�����b��eW���SCRj�憐l����(�@��`]~ ŧt�ĉv���씥0�H�U\�.tZ��g�l甗	P����́�$�`p���Ź�f}O�lT������-r�l��GR"&��?G��K�g�QNw&Nz�뼷���ɷz'�_F��V!�â>�����j�q�w��yXU��
�J|羮��yӋ��D�����A'�����Ay�d�6��Ă$�!�F3�b���$p�z#o�]�n�j�S���K��6��8c �ب�/��w9�-�sM5��>�K�!a/���s����/���Eِ�>�Ӂ�9ԭ���܎��8���� ��[�>(�.2���-E�{��梒O��h��f:��b�3$�9���q�n���s�e��p�G[�ܾ�fi�ˁ�Q����	ܿ��l)��)�R�ȶ�gy�x֖��x���?q(�X]�1&�9V?��j��0���r���F�?��� |;�P,y~U�	���:A#�vd�)"8�ێ�
Ck�i6ݮO�;8~/��FVUXO����w��~����m��u���"���<B��G{�3S��}	�[m���e�[[�>�Х�ܑ��ըP�s__H��q����N=�\+�F�jh��9�+LZq�p�IY�)���gf�F�qZ�7�������V�g����4�I���4�蟲��%y����D�/��[<G���e�9���W�g"~^$�ڕB��;Ji?A+�p=��+�e��'�C����Pf/X�.�&��Y�(�ڴ��3��ơq��ZM �&���y�	*CǼ����41`3u�r��G�J\��q�t^�+�Ȭ�y�i�:TҠ@.hy��W�\���q� �c�V���9w�ǫ��� ߃6G tpT�V���*h�N�`CZ'�;~���]#�aˌ��F��9�>��c���]�џ��{T��Ψ���t�v���;a���z�:��thL�$fϫf�'1b��� �o-D�O8[�
����gs|�fX�C�X�	L�kY_9�o<
N6$0�%��#Q�z"�>U�b@| ��'+�f�Px矩�la�!�|�P�xj'�֖�@��u������Վ��9(�%���=��v��mUAs�8PG�r,P���Y.�g���7�=�4��!wmY�:~T	mKK�g���"�$C��p�ez��HA�@1mB}\��E�3�������t`�����`�N�*ʞis-���}�W�7I�o��n{�S��\�Ap�и��9/��jҊ~-��_ɵ�P���.r �6��0��V�3~�����cF�?��^ʳ]i��X�nQ>����@D�3��5r
���VO���AꚔ����ʤ��X6H[ "}<E���wj4,����Q,�=3N��Zy�U�(k��<g�s���8�'i��(/�����A���4Fa�=C���0��"w�/0�N*_϶���c�h���U��B��E?'0��8�J1)J��l�R���}z?����R��ı}��t��(@.�e7��$�O��l�[_@�5��>2�����<�����}w1��<&1�y�|S�m��N�5��Qp�S �7����ڭӏ4���n�{��RZȂ��%|T�:m�E����{��^�F*�����D�	�(����ܔX=������R9#v��F��Gi�d¡2z � Q�I{^|�o79�mn{iT�j_�t\{ԇ<N�Wi��6y�4���񩐳�h9��l�t�%N~B�<wjܻy�͹��s"��D̢��Si����`���hCM�!�5D��ɨ;�q�;��H�0�p`z|��g �;��2Ӄ��nA�o��,��|P��f�{^�9��1LO�\��K����v��OOGW��y(,o�^^W%=ݳ�ocK��*>d����4�s�Ԑ��O�r؛�u��)n86���0V�/�i����CI��2�4K�G���R�j�(A�}0cƠTO���C����ֶ��V�1꟏��֧p�S�}�2�O�#�5d{c��@�p�lQ}��끠��sPS0:���—�Miu�]�<���x���Φ^�f�!.�������[i�g��hQX3��$���P�ySL�Ŧ����O��ӈ�)%iq�P�zkˑطR�']_쬳�)V┩e�1<�8�D�����L=���2G��5;XL�p�,�ٚ����C	r|��`����̭OE���6Y��T��i2U��d�X�����a	����kGrݮ��R� y�����U6�1H/ ʳ�y�(��.n��C�R�SϸV�N4�о�Ü��d�4S��]<J.�+�$π\Q��L�'�O ��߮��]�d��~�UN�(�w�PE�;�I���\��˄H�.#�q�����g�O�d�^9���`Uv�������蹇���|*ρdju2�����o��M�ͷ�h�O�6+����x�Ͻ�#y1Ph�"��ѓ.E��-�1�拦+�T�H�4r*,��u��%��� |/�HsVo7�s��^��$Zo(��������=	�ӮZ� �T�.���^�J����
^��z�0�HO෧z_=���9$�ܩ\�[B,�0��=���)M3qo+ 8� ��jŞ���PmZ��GeW�.���j.�3_
�N�$��g�EJS$���k܆>AE��\�Q���L%{��u�1��d�؃�b�O���b*�l�dp,C�lXƔ������fc�D3���ٽ�\h44S$5�L�,�1"����8:C��,w��<�E�g{����˪��:��u�[�V�!|v�h�O���U�F]*���{��� ~N!Op)�~�!`q�
�+b��v�1���4M��}M����M�J�,U����T��EѲ��ʀ�t�������s����h)��S�K&�r�Ţ�ly[���|+}h6B�Ӡ�}>�ם_S«)`c�l��MR��/OF���7���j�]7f�/�z������>�kJR��dw��'����$���%¸�ţ�
���4*=�Kte����]�KHc�Lx�Q��������e�`�"Β���D�#A:Oz! �u���i�礗勈%�5�a�R��d21r�}Z�a���@��>�p��cP���]fD9��o�<|,ہ-��;�?�C>s!����Ӟ�j���9�g�~[9U3�U�R/��"��'��P[}X4�
�l�Zנʈ[���8)K]%��\�-��e��.3U{d}���d���94�����!������-+�p���&���^���"O5'���[��*Zl�{�	)�%,��A��%��HT07N��@�K3T���0��
��wD8�>����H'9�������V�e����Gq9�jkZ"�<̛֧$Tn(�
}�락vF,��-��#�of��k`n�T�A�qL�U,�/5[*���˳���R����V}��/-Dնh<���(�7��FPp�^���*��\�iÆ����f�Ŭi�P�\��POn$��-�����S��Ԉ���2&��u�Ug[�n�!�̾R��w�D<_1wyX�X�4��S���>~���a��7�XV;���v
�+�Rԑ"��uz�oo�U#�Ֆ$t��[Y`bE����\��j�.x�D^S2\��Ɂn��e�˥54��Gd^�	�7���P�Ӝ �h$YP΢a�#��.���R���P�@6�r8�S?m���yy!b���b�A�Y�
t��/J�	�qˍ�-��
�C?�فapYB')�G	�]��#�_R��b�I��J]۱ф�",ь�6�z�o�=VN;J��W��6�D"����mR�V�d�=�/㟲4LҨ���$:�tE�8f�⣕�>���3�kĐ'�z�>�vBG���V�q/���3!<��1�N,}���t�P$8�����Vm; ���Eb�-�#3�5(�28W
������D�l�q��i��_+t��U�����ҧ(Ҫf�5ķ��ǅ� Y��2-��h�	:h8��{���y�95b(�#	)�L~f���۵�Z��l�-�Rf�\{�=��l[I�*~�������E�cë�`�x�!)�=�F�۰�[�R�c�PfF@zbV�4��醬cZՠ�״����Z��)�1����>�"���2�I�T<Q����[q*�f��*~���W���gGs�c ~����/��� H3�5��P5�( �[TGZ@-�iʍ7��V0�PH�n!޶���vo?���=i�i��3}#��q�3��U��x���E��e{k�$��M|!,�6��PEL�a�5  �ݯ�����en1e)��F�㰛j�kĬM�a�%��(��We��2b_10z�n87�s�9Z����V�#����g��@�"}����'������w � A��_�:�^�=��1���@��h,82���%�$�n�V��P!"=�޾𫶥������:�g�J��
^�_ļE�Aq̰b8rF�J��Dᒨ�	�{ҭ��vZ̆h�<����Qр<�UHt޾&|�����Grw+ɠ+�ﾴ��,=_� )Q���� ѧ�mM�m��!�K��ΐ�Τ���$R{������y����%�	��n��-��Q��fHd�a�������=;������`<烳��d�������ދ�^�T#"(p+s�e)��ڢ���砢wRH�K��*?�u_/ׄC8a���r[n�UL)�d���@��zZl)h $l�m��߁��W��'_$]mۜ$6-�`�S*�Ha��e�����9�,����0k"�����1��_D���z2Iw$|����������H�9`*�'Y�U�0̈�bjT�E0,M�r�G� ����R!+r����@(>f3�	mݖ�F�a��G`j$h�ab$>� `nYˊ��.^˙b�qi�/���-�k�ZtQ2�q���l�{�t���B\�z�8���~�KwN�.�ǁ�Z+�%�����c͂O0��$ғ���ܿ6S �;���b����%��Eh'�5�lN���0蕶�#ʆ{���uwu����Tf��o�C)����4���b0�_)Ǻ��D�0�ugG��~���c��S��bJk@�T��������Yv�p�㍛,���M	A�2S����ųQy�=�u=�TIk��pҫ3(XZG���E4�
����^	dX�%����*�A��t�h�EJG�����L���O×z;�$X��L_T&�˦���}���=���}X��L~N,:l��$���hH_�tIxIX4�� ݘ2MD��XI��,OA�(����ГM䚊�R/�Х��{����Aw��!��,��ג���AN����o-��h�5Z��];�?x���Y��l�^Ӭ��9�l��;��J`;(��a+e�d��iT؉��PZu!S> ���z(m"��^ʽ�O�_�B�������˱�]2�V��=��H2q��Y��?���J�"������Hm�a	���FNS�|�\h�?�3fBv�iI7��ŋ�4�g��]N&�5��y��#�q\�莀��1_�q�@�m��eG\��V�xp$�	x�%���Q3�"�y�*V��xW�_"��P��{��w���޵(��������)�!��D��2�s��|1m�ɨ���z(΂�Da�-?+#N�����"�͑D�O�N�͎B�Q��Ě�d��W�'~����o T��F�A��͋UN�ߒ�|buqb�e��3 �C�k60�# �a��o���xE�y�u9��f��y� A���L��2[���1�
��($�-嶆�
�5)�H�)��<d/I���c��'3�^��h!�?�Yʎ��.�uHK�v?5ݱ����56��L?M��_��݆�.ݜ����MB�N+��.�TU7����8���Gj!TI8�x�z��&P�t� �<TkB�*#3�����
oV?w*�p�e��N*���<��{�7�1��=�����ܶ;֓�jWxFG���9棌&f�(�p�Lg���0�?�J�JIw���(S�����l{Muh��a��� SB��^�W�&w��� K(��v�x��%1�� G$�U�2�C��$#�j��1�!Vyet�����G�S>���]J�Rϭꁿ#���TB�A�(q.I�=1�KG:pW�~�h��tW,×��K`6K���f9���'������J��o�e�am�k����1�۞"�{�	��-�:1��5�)�1@��РE�W��Ŗ���Q����/n.�&K��+ /���9��W����S���Pe����ct��eap�#7�@�r$�eЧ+�q�K݃�Z��;p̝gZ���QY���U�(��+e�K�>�:�L�u�fl��L��k�/vs7��$7H�Z���������
���|l�l�5�� %�-�j���E�*͆��`�ߍ
�%�^�N.��7wGO�YVn���.�ײ/��NyE�9JR�6�V��)�},�`��8�fq6s
��qD��8,~#�1�Z�O����bXY�n?	Z�(�?�
G[�5�K�k,�ӪV��3����h~�ſk*˽��!y5VrP��i��D/��\J4Ǥ�j�d�'�J
�Gb7��@9�O��F<u��g0�ò��-_�+��$�tJK����(Po�����vCA*�_$ �k�_HO�������Ḫ�F|�]�,�[��DO VW"m�<ѽh�w9���8P�)wD����ē:�*<z���K��YcM���e�N������r��\5"&�ĝ~eF*����48w�M�
�E�`���l<7��Єe��*��h'_b��s�'��%p�I-���U�!���ˈ��NŻ�f�m�m�#��e%p��d�ю���}���<N,�>��R�F�����rN�u�˙��<�f�ո7l����7O5��	�Q hwtB4�8p��A��qM
��OJi���$�r����w9�$��Q`R���б����U�w���- 1��ʺ�ώ��t�I�WS��g�9N�D�ԙ�Ĵ%�F�*MZ@ML@zd�,�S�7��F�|�F�&L@RMՑ�;M�>2��s��� ��p\[�=�D[mqMX�J�����\����3C��q>�ú�j XE��!_�&i����H���`�-l�8����Q�'x�Vǡ8��o 	�zw���C̖tQН������1�b���Hk-�ϖq��c�bh5�B��p��1^�������dÒ!���ȅ߈���x%`Yp�;���_�NV*��^a�؆t����O#���n�y=���~�ļW��3����(b!K�,KK��j�~�ӹ��X��:{��WcO��V$�[��Ǭ�V;i��ܥ���XIlPE#_�-�����S�^a>(�i������)��?���X�t�b�y���M�̱��C�!P*�ËU�x�l�
gx`&.4�-eqgۯ=��P���N��JS�"�\V��	WT������͵�������R���-QnW���)��-v�_��xV�4�A��ܸ�$�)��#wH��_k��=�-�G��@���NЬ�d����j�)������b�S���q�~1m
Q��^��3�&}�B�Z���y����bp�N���)���N֞t�&g�N�qI���z�~η&/���|ͦrC�?�b|�W����o� +�_�	��^�Oй옔b�Q[Ā����uq�V�����s�6�EOb�輠�)6V}?Fh ` ����c�	q�f�8�i��jRu4�}U+հ��Y�.�'�QƸ�D��e ߊ�����e(:�=B3p���ѣx���3�%�Z���M��DV�]�]���y�uS�o���͗�:��xg#C����]A�B����J����;#���G���$����V��LB�J��<�]t
4_�HG�LEӑDEW�*�Z����먋$�e-��_�Y�[a���AG��u��C�����EP,��Yݹe�_�Z?�b<D�w���Җ2���>e��Џ�<��)��7 T^nHTpԏsA��IQ`qjJ����G�S���˓�ꌢ��.�5�{D�t���;J�RE�p��ں�g�סF�kk�X���H_ݻ�
��u�\��ڌ����8��iS_�o�����|2{Cڭ�"Z��.7꾙��o=�Nح��ܒ�iQ����g�]�:/�ĉy�Q+�Tܒ��m�*��q���0��3t�-A{�f���ei����H��)Ϭ�A=�s}�l����e�A�k:��4`h�>�8A:X��$r��~a�R�N����Q}��s��3�}��v��=<�2|U���/DS���b3�	�%К|=���x����_v((ܗb�.��<'T��`o��*�s ��Z��q�/蓫k!I��]�^�|�ޣ��W��m���1��^+�羿��Q�Y��Iaٻ�Ȫ4��ڽ��=WK�Uj.t�l`����J��/�ɜ�svʏ�B����Ut� ��R-I�������ly�qk�\Ӊu�԰q��q8ɨ��kC
�/7�a�T�;��������֋c�yZ9Zn������	��Y_0��t����b1�'��D���FɔR�,�<&��Â����s��^ �9�ɖ��8�[���B�0_xaOF�M��s�	[��2`8�킕<�#��B9b�8�ݍ�-Nަ�J�ᔾN��n�~^�A`�[�Ak�'A��l��4����º���dU���02�Lf/(�ʹ�X�xK/���w��QO�*�S(�}�9�3�<H9�8��%L�t�x�y��I�ga�C5V�s8��D���dJ;YnO�e&�"����!�N\�
�;�y�[C��)��@.)� ��S�8�I�p0^VLR�Y��,2�')�T��s���V�<���Y���-i!G!"����0�F��z�#��b���[���2�xw�՛؈��ظ�
���9V8�>�=b=~S�(w�`�����9�l�8��ܬ�@�J�T���ЋqH;�_W��Y�-�D�Y9����rn���M�1]@6�h�3j��9�Y$6ZΓģ�唛��p�uF��5�\BKg��(��i�Pz��.�[��mZ���ts�z��9?%>-�OTZ��>c!��A}R1<�>}�OL�{�p�_
���gUՂ��W�����$�}y�zȹ����Q������f�������z�zB��P�IWT������Z3�݈��ɑ��٢���e\R~wi��L��k��#�,3�tSev��ܱ��$0�^Rl>��P������<��L���
��Z6j�W� z'��A�+U��� �_�b���V�"�Q���k޿���U��=5ۿׁGa'��6^N���qh�E�W=q�1�Ln�I,��)��x`�]�"��F����F��y����E6
H�)�%��0�r�@���%����D��w�R?�F�QV)��c��b��i�S�ǥ@�h�Rvn1d�ڎ>��"��?��&�`-G&e����4�N�#OS�D7�-�Ʊ�[�b�Zg�;?������k��zdO�4"���/��Η�8�-�	�,aDڼ#B��"?@���O�6x��mXJ���JM��:�LJ`O�oFB\2���ؔ��}�3��J����/��eH�viReWb�Ţ���^�j"8� �jK��� q(���`OY!��'z�˹tT����l*k��-%�L�q����^Jۇ睟���R���? �yAV�>��=�����@sFH�J�g[Xr�(_�+�ʡ��/ݑ��u�kLB�KKJ`Z�S ���,c���=�=�*D��c�xN�Xvr�)n[xq��H �uá>�X��@�_��_��b"��P:�s?����ώ92�Ʉ�M�������s��I'�!}�~��"u���֑u�p�4�E�����-�WT��<)����K���"h�i����vH���5������<�H*�.T|�v�OњR�#���	_���~�����]�����jX)']�\�V@Q�G.����tu$5�CR%�[iyۀ���ll�<����t�4������
�|㭍.S�JZ���w�{�Q�!Z��nBCɷv����D]T�d*䆉�Lg��x�x�7L�V�#.$�f\��״;�\s3Z��r��������]�z��{S\@>����ٿ՗��8Z[��$� �+8�Txw��)�Cr��#�ͯ�����c�X[JUA�z�\��4.A���:.yn�Wv�j���@���S���3Gw#Tju6�7����d�9'�d���#�a�6�l�)pᨉ��6X��\^|�2MN֊M�]2�5���9�� �����1JS�d.K��)S@� ��h���S|��
iC>�T�{iI�*��%��ƶ>��7-oQƖ��7�Ux��,�]�k"~��ឈP��	Ϥ/����'��=�|3�e�:�[o �g� �S�Սɩ���ר�6���ms!Q�����S����z����*�w���S)��1�ȩ�D�䑍�@�׆�~�vNk�P��r�P�g�l"�R%��;�#�T�JaFֺZ4���d��Q��9�:m l8�5شȎ_��ܾ��c(t�_tA�o]\��~\��-/A�+G��<�o �.N�@��D�w�q�'�H|'y�rk�@$��{�*&�v��L��oi� *��+��'�p�=�E�:�&����2'�޷��:X-�NLkX��D�*�Ղ!�����֠�K�ag��v1����μ�l&��^QP��J�*z��݂��:���\�ۗI��"C��Z���q��חÙh�s�|��Ƈ?�*���A�������`��]I�ݖ$D�iq�7���b��mQ|c5��V���C �EC���G����-�u�������C��8������b#�>�s}�3u��ԩ�*ȶK���;�/}x�2E`iY��r�2Q�Q@��%٥������s"������^������| �s?���������C~�W��Kfӹt
�, q ��H��(t�+��H�V��4>����zMFږ���v����[[GCx	��!�?��x�=~m6͕�cy�I!���2�q����z@G����lj�=RV�e����58޴�9�C�|k,�9�'��T�m�w�w^�O����@������Q��l!������l$��B��ȯ ]�q/8 ���u�+�S3�bcj ��06��5 tE�g+��Wĉb{�T���gZ�����~�Q<_���D��X�@�;� �[���"�CI'�I�H��w~F����9�Ah���c�w��Ψ�����z ���ٜ���#�' +Ʈ�1��{�Ema.�1Z��5�BJ���H� �u�L#_�a��d[M(�s�݂@��%�x�&C��X�h^��ؓٸ�yI?�t3�L�!���7T�b�C7۟�R�ҿ$7�l�P��`G��� 10�ڥ ��:��sw�G�Ǣ������yiZq �#b�]R�@�w� �*ܙ0!z޲�� �S���u���'�K�������\JH��ڿ:Б�D�kX,���&�1��w*�kF���V�+�O�A�F��H&�A����2q8c�����[O�����
��WG4��w�Lë��;Do���G�&�4Ӓ�×������]UO�Ɨ7��%�y����B[� N�$�>���LF���d�<��ھ	�Iog:��Q���K�*9��L�}����$�r�L��(�h��#k�G1����W ]=P�@���6x�fqWRf#�%o��"