��/  ,�8Df�E���f��Tj��Q�ˑV��)�ܜ� ?�`k�(�:pc�ֱ&�T��E� �#�ءO�����I_�z��Q�7��T�)�!i��ힱ�fT0W ��g�����y@����Y�Z�����?U��qӘ�Q(G�V�/_e������}�>!B,$^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK ḁ֤cGG�	�L�6�utB#W>�4���ո�����19v~��}����	?å~@ ��ŉP(��eS)N-B배������Q�>h?�(ɰ�Z�yH��[A_}n�٤X����@�BW� z���l̰T�m7�"lZ�GP����|���tQ�T�����&"(*j)aC�A�C�U���!���.��a�s�l�E��y�?�;�k9t��SS��3|g��NT7Xty���=b=%��[ܟ�>�V
�5��)��T�8�P�/P��2���2J������hG�v/�:%a�v��Ȣ�:7��7|�fk!,�i�Qg�!o=� ���7�3���A�l��M�\{�2���Ln���ͦ�UU~�M�1��E<��Ԛ���~�.aǒ�}w0ؒSv��(nk6^c���-IKć�]6|9@b�Vr���_{^t�&��T@S��>҇��z�w�3�7��^R�x^c3�������y�nԂ�#'�=��G��5�!�]��%%�Z>��M5��_������7	�n ��"2>�4J@|֌_���4�%pa���Hb��4�@��UK��^uGZ3�̾�e����W����'nl#&3FNP#�a�'{�'�ZF�S���ɤ45nG�i�R����k��=獴��i;����x�>��ـP�9�`�B]�c��ș0���77���8�ƫ��V��'E@��>n86]�%u�����lj�!'���/��-�ߨ�gv��J�*`��$O?����0�$Z1z�֋�h8��U�vK���Y���PQd=j-�Le̭:+I�!_IȌ~��=˘�(�ؓ�X�[�z�p�A��`s�^R(���w�5)6y~R�,��;ջYsf����.�f��`4����{�O]��!�qϫ�F*_Br}�h������97u�QC�������O�jr8'�����T�>U�~`Yۊ�V� h�E�V4t��_�M&��r���r�K�8Qy������cg�oy���s�gi�#����0�#����G�]ث=�R����������=�=&73,��~�+j0u}9�h5a^}	;�:�@��������X5}�\$�v
	5�N���c���� �<P�.ޱ  �4����x�m�@)|��@��9�e�c��S�6��Ϲ)t��~�W��D������aҠpu��;�krc���4�[��Xvk�/�5Iv�[��iB�O \#�R���Ӂ� ��p��H��Z(�{b�7�.�5�]�XJg�;7A,��р��ߣ�C�n�����Dӛe$��|?ۿK�?j
L�+��[�Ɯ���FS��Up��JZ�&���\L���(��uKB�H#�7��>Z�L�Wq%O�eB��S/��˶,�?2%�hED���rY�P�IS���}UK�9t�w����$�@�s��j�1���ަ��;��9ц �����Ǽ�sN�zT$"��n��'q��pٌt����΁���|i8jI"�q ��wuKCfg��D�` �fg����א���[��7+1�T���;���|}k����ַ�tK�C��44i���7VZ����r�r��k�]a�jgd�D��b@���˜�\����z
%a2E���Q�F)W4b	v��g	&j��ɮ!���&�W��3`㝰8�)i��C������5����z�+�^�1x�ZC������x�q�m�{Ԫ
�uo�T�cI�x	��,�+5��p	0�4]~��� g����.W~�9̧\�r}�����;̴�(1K��m��<_J�e�O��#<z���L�қ��C�A��]ԑ,�1��)x  =�W��w�����=bs
��ȍB?!��ι�6��L�=ɢ�e�)j��|��������X2����6�C_���a��hi�֘ Q"C+�B�Q,��ua�zd74TYt�fQ�����}�찴`���ŀx��ɑ�C>f�ݝꠂ,�Uů��U��i����1�Z���=6�������	�n!+�`��r��	��m���u��:c��[aR����5�_�d"�ޏ��?�4�,�v�U�5�e�怌1���B�Z�mhw��hv���rj����[�\�x�ٳ�UA��� eF�N��0�ޓ�~�-��ހ���"�2�K���U���@�AA�-���h��S#�A�s�	Cjn���#VJ[>�9.Y��6���g�> U����W�uN�Ԡ����||���aW��8;�@���;v�?���C���O��s�UI�"Y��B=#T*s�,5��YY�HJ0�[N�cˊ�fS(��N�1���j���ݭ. ��q�Ք�H��4�cVvX{�B(�B~
�},G���w� f�!d��� ٓ�̥�Mj�qV��`T����-�z���p
�Y��4]W���\$L2(9f� r������yIL!��ʹ%��pa�s��]KY,�Q-�@�i���}b��|��Ǘ�����|6o�� 2'T�b�e1�(���b;)���yGjL����4�S��$��.=r�"-gZ%�G�.���r4\%(|I��!=i��r�]����4��:8��Ј�*ɆS­�`��o5Ϯ<�/�V�,�[���������6������Y9�q(�)��_P0~��w���-��2�\�$%v �'���)���Ĕ�Ĕ��%w"�s�m�uўy��@�Kl'���[��_���&-�ٰ�ڙ�v$��m��SAGo���������<�?�D>�O�u��"&�O ��8ʜp�|�G��YH,�w>�#"b[=9�0{h�%T��\�a��fi;�W��Άy�֮l�ߑ����P�X�}N��_�4]8'm��8�eZ(�N�QxJH #J�h�C�{�1L�ڦ�0,�R	�h����I{f�+��/�`�\/�����<������ �8{"��:� ���~l>�5e���_��џ����]��D��^����%2y/��ac^��q���
5bL36�f�����8�.�W�8٘x�����Ü��F�(���O>bT��^�����,w�Nib����E!aL��h= ���Z�5IJ���>άԍ~]�R�ib`׾E�z+6y����3:0�L�(ђ'T��!�]�3R��r�*�T�8[V��ms�%��8;s�2����n������22+�y.Q�V1��jܫ�f׍��u�k�1���lM'A涕A3@�ޖ��<[P����s�r�0�po�Њ,�^�yD�˦�ɣg�u�<e�󘌚��R{�S��?��
��cfJ�x �SY����R���vk\l{7T�
Uf�j��.���Rk���߻�a_q}Q��T~-��z�9�J�����q#��0$�.�C�N5�a����+m8�~���%�	V+�ݦ��g�/�xt��g�Z<ŋ�Ѓ";�o_�$�A��L]��C"B��*�r�x�N�32��j%</w���?��	�v.�o�SDL�������g9��ž�I���"S�i>cr 
���|��K�d�UT�������^M1K����uy"� Nd��^��	�}�U��7iC�K����f��1s'�(��O�kk�=�Oش#�È4Q��ie�P�D��4|�wNB9H���Z��5f(�W��kL�����i��t6(;�:-���%�Q۴ݜ�]��j7u�2�yc�Nʬ��%	�*W�t ϸ��u�6Ę��vUS冏�F�$Mq�.Y.��;�0�VYB_�cdQQ�u�Zr�,t�ě��6�Õ.)D����'N��18����w�[�u�~�º�j�@s��a�g�,du�#���|#�ōa��Jj;�>��9U_�6&U��盒���˘�b�u�U��;�r�lI�!թ��eکFt��r������qg�9�g(�J:�յ�����oY��z��j�k4���xHdcYcW����T���Ø=���5H9���~�,� I�0�03)�[6���C�d��=�چ0�$�q3�t��D���d��#،��M�KK�6Y_P`���5M��A�Y��F�|C����r��h�W�7Y�c���3~�Q�Ŝ�O��)�R������Ύq֦o���!][Q�<(t�}J��%(y����v@"6wN:�?�ŜN��!�øn��zMU6��`��r�����=/A$���|O;�Z��!��u;LS�ZP[���ȕ3h��(���w�!����g%+�Y�3Պ�4A�ͣş�#�{��Ǡ��)@V�T�8P�#Q�z:N�7�	Z�� ������ �����=g&���p9܏��O6����>#Ŧ� �P;q�N�h:+i�ݖ�����;<�T���&���g�� �!=��b�c�	�H��'ݑ�ii���_�@��_%38�FC�/�z������r�Lv{���
Q�l`I��,��i��[�m|����I�)FH7���Y�h��Z���Y_m{A��Sj�C��.�������%e���Nĉ�n�g���n)L�����Z�jF�D���F�w�������Z��a-7��x'���Pg�F���g�=�o�͈\�?`�N���{�i�<R�����o��J/���Q���Y���s�ibHޕ�h�t6(����ޯ��1����I�)���F���'��T}�'�:�A��گ�
��������u>�*�'#�MT��j��#�@�W���{�f�Ք��Kb��qU���HR���;/�����0@P�c��3�6����em�bW�h6��u +ҍZY���i����B;6����<&�_2;
��
�����h�f��$Z܉�s�l%�[
w5z'OMe�״N�xa�U�yȋ�B,	�"���ӈz}��ً���j:M��ҧ�Ҋˡ�΃���~�Q�#:�y%����G���3�S/�2
o �qW��<W�E�Z��tV�#�H�/.JB#I���'/B�'�A2˄0�W�?meTP�9�u��ӏ㚐��<�J�y/|b�Z��@��Y��? ���+�O��h;�m��!�S��{*4�%k?x#�B��(�U~���6��´{�s̨��BE82����z�Kz5�#��P���䰜�D�~H���y��+�y�����tѩF�������8��..��E;����U���8�4��Wz	l��+�8�]����l[�mLT��ݬ8���T��u�4�3R��J;im�}v��o?�JҮbr��Hb�7P~�`��"E��xc6�ԯ�p�ʶ�/TZ<��*x}Gĸk/��X����n~�9`ղ9�]�IO>40_�s�%�߯5^�A��*�Ht�t/9e᣻}wq�P�7�4���|ڎ��V�M�«�X"��_V��#s�(w�Ge�f�R$����) sG��é�=b�GM��:y�Cs�F���5�]�-�.����`<�1�q̃? �����u��;2��}-�������t���ole5��l����|'��`6>o.E�q?d��})��?����jP=��6�&\va��A�d7tV�0ɜ�D]
P�J*�r�U�a�m�H+P�n2�W��⌶dt	!���\cw���a�і3|�+ 3�~��H\�^�{���A7�U�������T��a���*�ة���w�qh�8�R[�I`�N��F@O������?u#����?R���K� ������e��@F��]����r9L'��d}nh�#k4���(��x���:J���Ym �f��k��D'w�X�"��ӯ�dݲ 3`��1x.� a�F��l��p��x��s#����j,O�GC��b�v��6�Gޮ�'�/���ɂg���3��/��ckY��Hf<��S���@zK8��?HAތ:�N�x�(pu/�{�/A�ױ��;����FL2O������G=F4L�
�1$�.��4ƃ�m�@э!3t��|���vV��Ƙa��I���&I(S+j��S~�@�ǖ�0E���P�J�f�iы*�o�8n�C���}l���yF�����&D�J��*��V����_��xf/��N6C�����2�"NsE2?��O���ޝ)vr�קV�� w�Rs����C =+nV�_$����$��E��V$���O���a&(CK�V���[9aı�ߢOuy)�9��B�}�jIp��k)��L3k��!��ט�lgہV�
<q����Y"�7\{�R$��t�f���k��*���z�E щY����ُ��l����>Ҫ	e��}TZ뼍�(�]狶=.�?Dh7� �KJj�#�v����*��} �bYuT]�~��zj����ةQ���K�D��	"~_����.MK6E�;�A�[N�=ȝ7o
�Z����n�ھ�Rcn+?hVm��!�T��љ�#��?�UuE�6�\���}����ʃAlJ�f���bVW�Չ�����6�J�l���P�禨��y��a%�* �T��~&�0t�?��w<�]�~�?�0����������! _}3���!�f��e2�Qa'��Fx����������=��_����r�C��V���9����q�W���'��ϑڮ�"�=��ы��M6�3�[k�m�])����R�B�;h|�$��"�5P����R� ��T�k��
����g&���,�����މ��{�bf���5�Dv�%� ���=�k^S/,1�,5�	���.#{�4�Ŀ+�F�v�$6>y���΁�Οq�^1>�����}cƶx���(j�3u�¥1�8�5�HOz\��L}t~e}]�^����B�Y�҅����tR�ʞ���ua�[�H9eZ�-R�9T��H�u��gO��56T��S�w��w᛻�c��B��[��Va B%���!��豠�;�ϐ�|�̰jY���{�u���q%�2X�=��?*Q�L���ro������!�榡$�y��+G���e�b������r����1	е&Я�g�-RL���s����s��Fu����tx�qLYVBc�#K(�����*n�w�|�I�� r���&?-�o�G9.}��/&uՒ� ǚ�H�G��]h���9�q�iFW�V^Ճ�,2a}�.���HGK��D�l�n�6K� H�o��;I�#�����>��%��ݍ'��Q	�紫M[~�TH�T�~�I�}+�rĀ5	��̼l�y��I��8��	q|Xt^6�p����%,G�ȳ}�'�;�ciP&V�.�� ���5�,�=��[��Q�4���| ��}��Yr�0R��1AB��cd���?�	�"�4�ך�r,��&�
�"�g�;꬀��ǒLUQ�mJ/ rE��-�Y��c-�!+z��M�7�Y�J�VF�?��%j�t����K��U�m4�jc���?�lp5��l��Ж����u�p��J߶�֖����<tf����� ���$2\��6�_+�Vު��M�r�X&Mo�(\��J(C�]{i���[�Ï-�9k�BU�,{#���b�����	�����Kŷ��(e<j&�S��8S��4YuO���|@��46�������Z�0{��#�J�;T��H9����� 1�r�ٿ���H�;2va0p�L��GG��ie���1Oč������'L�PXQo�j�����/a���V/��H郪*�71l���i�����G��3�X|��с��h�*��|z�����z�{�Y1��0E�%����e�-NC�)ϯ�9�樑�O�G~��2D�<H	o��05�������s/�Ȫ��+p18B�u�����X���"�%�j��8��M�	w�g۹�M>긓 ���%mV 5�>YG�잋p��<�+�����9�sA'� �֮kF���֬��:Ok���,���d��6Z*>^2��*
�ȗƳc��-�� �U��l��b���E�w1�^R���e)s��dyzg�"/F|f�[UapG�@�MM1�^64��֡��}xˍ�~ŋ��y�ǿh�ܵ	TK�m��V�4�g7-�gp���"�@�ϝ.K����/�_	܇�4?HA�d�r{��,D�SR��p|�yp3�|R�Z���lM��JQ3Ae���0ҭP�J�T�W�_q� ���Y�c9ǕVf���XX6ZѤm�u	)hvc(&tf�	��j��""�V��4pV�?/��=�'*�#H�[��P~�('-�0�.�:��_g�O�<�-WC��DS0��� �\�C�.���/�M�{
*�m͓���%2��>��d����������9�Y�چ}7\~��f���w��?���g�L�d
�:�d���G�+V+s�?T���Rr�e�3[��f\G��|w�����/6¿.,����1�;����(���j����)�����(��S*�Vl�����Մo���{s�k��CUo������~��}�*G�km�r��-����n5.�qH7������bj��Qs�qr�y>[��r�UT	f�%���r�/N������h��)��0�s�U��j4�k���ӛ��g�H����g��(�������Q#�^���ax >>���Q��?G���>q��5iנ�{������'4�%� ��WG9G�U̲8���XG�jLtG\�K�M�T���4����V�,'���zp�d.a�5@9�B�9�W�(�ȯ ���r8��3�x�,��/y�ۈ���1�uQ���Gɇ�#�13�u�Se�� ��ǯ����-60��_�16׮ǀx�։" /�;fG���'{��Xq�������qU�l�������?��u�/;�٪�B��$h�Z[b��Q�y�9��٨-����1~��?��r���8 6H�7��s�W�By�i��K�x�.�6B�j�I�VW9�]�~�Z�8B���z��=�x&�U����99��ﶠG�l}�� �;����h�n����P
޲�^[E���3ܣ� �P�$mD��3�����R�h,��y/��9a�+�Q�^� jB'�7n;�U�)�	�uZL��"W�#�c��&T���5O����h��J��e�%f�%j'��}1)��	F��	�g��ȚD�Ӥ�D,)z��2t"tV�����q5,���OSp4*����vD��?$j�������9T��m�A?u�_-s@A٤ :�졁if���dz�ـ X��9��:&r�F׋��0С�ڳ��[5�R<�������-�u����r�3���¯im"�"�Uw����44e=�0V�� �IY�7��S�U��B]$f"�t0`���w��S�/B���a�],?y����H�?֯�3>�N�v6=Z%g�9"�Ƚ���� Z���l�W�:6�f�~� �@Ď�}nIM=��7������z�%�-��]�I�@D�"��$�p��3,	�Wj]:��3�����v�R��@W��Q6"�g��.�"��e�d� �;����9n��z>p�Ƅ�>^����6i�(q2�Uui�Jɩ9���qD��/�z;
��<��P9�,~��d^b!\00&u)NĄ(��� ��`���S��Q��X��H5;vF3��\
d�b�NE����܈6��n�C��f1$�.�/��z��w�d���J���玃>��P5�-�SlD��Z���%�3����T��Bi��{� �&�b䂌����(XO�h|����$L�N��J�����?S���:��K�Γ�b��Q�)�^�{�_P�����q`�V4zUGb�|ٿ{�@���הJΪ�?�/5�'��9Z�v�A.����x�0��#�SW�z�������XI�:K(�7�i�M�i��ms16	�W��8K�E�M� ֖�M�CJ�ێ�)r*�4��V1�
<Ǝ��_�8;���S�8����.���:m~rg;oj^�R@�'���%t�fa�������l5�F�9� Xh`��6���|	|���XQ��Gh�]�uZ�Ū)B�Q[
�.�E�hZj�mgd)�E�[�ȲD��!�8��Z�B2'�K؄���@a�MxE�`Dy�(h���dKSޟ���G/PM��6�~���s�CN(,���	?����wh/����=���1r7#�Ya��C���y�|HR�tfl��'���f�d:��MOm/p�О�f�X,V2���	)`j@{�u�_,�X�rbUa�6�1����X�#N�]�����{�[kc�{R[���A���4]K��e=Qq��	6��Ml�(�;�����<�YTX��|�������q����zD����2�Y�4U�y[����B-����7蹥�,�
:!G!}I���I�=g��(L�N-�Q�ßI���g'2��R]��G� 44���4Jȉ	s���"�u޿kW��9A��5���o�5� ����@ǳ3�Jq�����>A�^V�s*����3�ۤ�Pz�'x�ᨼ~����1�����
D�U~�`�8�ʥm�ݣ)f���6�DVs�|��S�a����^�X��L�N�tl�-�� �$Kip�ۼ�@X�'�R���62�u���屹�jqJ���)r��8U�����8'��ŵS�Ygs���k.}􀌯����L/X��#�؃��U����СF�#RwF-��uC����^b�v���8��O�s�=�v���	�X:GL�i�������(cj�1D&Z ��4��9ފ��w��� ��`b]�oe�^�q���9<Həj�oki�ll7��\L��r�\���N�^i��f�iS7����o�}r�b���1\\��2*Y��1�0�R
�l���/��=G�r��n�6�	�[XBk��b$+SRl_�(	5���j��U�AU�>,���w�2%��Bt���V��E�iD<�:H�'���^.��1�ә�Pty�IxX72��@u��������fWz�-*��vn,Q�?��! ������Hk�Q����ҋ5���,5~E|׻#�f�l��������,?��O�K�gqB�F(2��ǘä[�@3#�w��� ���$�F�gXF�!]x����Q��khs�nZ��J�mE�9r���M�_n?�������Z~� Ƃ_�����T�n�3�b���8���Fb�!�-:C\
��4!���Ӛ̜�M�M��d���Q�k�E�m��f~A�:=�L��ze,u9�]hwKK���	Nj:�cw�#/D��ZP��8}J$�����ɪ:3Z�D�c�@�z`��s���k)d���ؙ��9Ϭͨc5���+E�S�Ɨ��:�8��݉Փ��a��Ok�Ó.�!+���v�d���wѸ�B@�B]�&U1t�"�V:���T���|��8�}ͩ�,6���#Qm#^s!�&�l�K ǫ��W� D��%�M�9��d��)1��'����� �N��u��h�.�(Ȥ[�\����tz�Y-<~`�	@�ہ�e��[������Kփ�N񸦯�!�������F��9>Lڢ�V�P)Lz�����i�d%��u'����^E2�a���*�_��w�p�����t�.H�5/�V�o��ҿ�O§4�[[�p����!8���&��ݏ���uB��U�@�
��4b�F��b����Tm����q����SS>c?9��M��}��,Ȩ�B��7	)H)�M|l}v��ew���\I��YRޔ-�S7��Ӆ0!��)�PQ�z�C�9Jo�m�cnznKgBT�3-K��)��|���b�� uG�^��Na�Nt��z�:\<�~�j�$�g��&a�j�6��|�N��N
D��Čo��6 ;-�,K閠a˱����k���(Md#�/B�4�C�B�}��;�TeH�� ��7�*��u�0���b[i^�p�I�ZQ�X���@e�0t�*��x}�?UB�P�
6�(�M��+���M#,��:;�ӫ��z&s*5�0(P��B	����8�����L���.�~��Nk_��BE��>41�L󸞗������h���t;��ӊ:�?.����m;����E������~�Y�Y���i4����Й�fs�����?R���{��˚��D�����JD�H����Ɛ�GFa��j.�J*u|�<�5,E�;Y��0�6���3V�l�>��v�S,�1�o�^k��c �t�C��:���F)��m���`�0���\�y��O���W]��B��%� ��-��3(�3�s�3~���;'R�W�r����q���v��?�*�G��_N	�ɇ�ݚ	��$�W8���~@y���p�4��W2R���x�w4n��*Rh�ԘASoh�v)t���D9�Z���:m<S>��ɳn�	e��i���f�;���x���\#��q�s��'D��3\���,��Rn&�0�_p��@ιx[��V�N$�8("���9 K��b
�g�X|�˳���_�'�"��o���χ�"]�8�S6�{���g�,ɲ�J
�i}8��z(���%�+���q��Q-���mI�mEzRX-9
-��dPT���I�L��=�v�<[��3tϋҫsl�
��SCc�P�D)UZm��~���ڠ#(�J���������h��rJ�,�m�)]�Ou�ʁ�iNN��*y'e鈛I�;Ւ���ك"�'3��uSլv���i!�hVIf<��ʉ�f�'��c(Ŝ�ɰ���
)����49|;�➨����q�NA��-XS���ST��D�wb���3�`�R���/���5.]��e�k;��]L�6]��`�F�/�gƺ��E�h+�N�!�3�-�H��v31��R+H@G8_��D��ݹ4��ŗ��"����7�ɭ��U$A�����I#�."�$fI�����D�1���/��[����u�C��LI��ӣ�� I�,Ym��m�s ���<�1��ʈ}���<�ˍ��D�-�M	���#i� CjD�a�rk:T��L�6�IyK?�������Nu1���Z�'>4�C��N��cU�>���"� #K�YZ;��&)-������a�O�ށ����ђ�m�.F��~�������B n[�8�%:�|��� ��:�hv����v1��LѾ	�{-��7����k�����[��ִ���w]��;�%^�s��Hǔ��i�˯�S-�Nx���s磼W�	���Jw�\���ֶG���}���H*���O]�Q?�i������|���E��.18���!��+V�=�A�W�:q���]�*�N
���2�p���n2������4U���:""�;e{y��q�'OU�Q�b$�a/Sx~68���[hP��"���j���~���k����.9����ڴ������"|h��ׂ����.޿N�:<4����TCC�K��`s� ��Ti,�ߐ��#Ɵ����\�L S��P�&며����6z1SG� �%�$^�zb.���k��q�"�?�U�|��+�V�xܝh�'>�m�k��!���WN������[a��l�	-��]��(t�:���r�Mʎle�#4��h�ȥ,v�����&��($��;����<��(m�m�+.���Q�FV�c�E�wث+���J��t5�{��gj�0��IC<sCgJ_�`�W����Ǔ�}�%���d��zO<e�I�����!y����>]jec�|a���xk�}����v&��hӆ�P��<��+��\����n��´4�r[��K�sZ��foF����B('Q}Z׊�Ju����S��ON���hb�����h��iI�x�K�t��M��[�c��ڝV̛�cvJwj��n�GKs�w�-ɮ��3ݪ����
<0~�G�a��z
��#��R'�ˋu�"x���c+����~h�� Uᰥ�;�����ǅ�n�hj�	:��@�A������[��7ຶi��FȎkS:F���Rᘦ=��G�p�ٚtW���,� �����xb����zg�B���e��bɆyU��Tl <,'�{m��=��Y��^��~�18�{����R�)�wy�'ѽw  � c6��6��jv��Zz��l;�C桭������I�\��{���S�{Ο��l4)�\kp��Q�8�A$���J�(l�_�	
�<pJ��� ���_��t[�� o�p�D7��^; �����7�>����D�,;wG�
}�òqnhZ� �E���D6�DR��w�Ξ�y�!�y ̔7ū2�� �; ��g�E�G��&.J��S?���;�8�MS����q`p�`�1�����р{R
��!�ج↩��$c�`;��}7�.�"Ԏq��E�V�>:��Cx����\�P �᪲aeU�}�?�{�Kb��ى�䐔?��8��[�}�w�tg}{8�>�QJ��iv�G��d��+ >"��96i�N�����Y6�3�M�w�Ͱ�Y gܴ9�`�e��&ݳ�w)ͯ Wh�'pl�ME/xئO��_���HAuBWY���؏7;��A�3\�{:���J���ը�|B��n���3��'����_�(*�[�yl��8r�3Ä��w�8w���^@����q��w�貓�ذ?��x.ͺ�񏣇D��"��Z���7|BFeL��QE.M�FP���ޕ>י���F7���`v>!��Q�s��T��T�P��8�����zYr%%65��N��$y��S�����H3�ׯt������k��Ү��8�!��Z�mN�ƌ\��֯���gc���
�T {թ�T97|Hg���_�I��ͷM��^V�sk\١�����W�A<ŢQ�=G���0�2n�op`����8}BdS`��SQ�a�ǰ�:���������[��@]��n��r�Q�}R���働�a�n^�&<���<�����G;vB�3!��W��<<6����wl#O������[NR��«�J�)��kњ,�e��݊�FA: '��M�`��*���-�t�8b栏�e'I>�k��*m]��F1�ר��k>�Gs�x�{+1���#���K͙�E�U��9XK�_V�"� �mg�a�@3�Mjsʬ��Q���3���]PnM�,q�_�NOMK��$)0�FCe@q�b���SUY�S��%B��[0TD��o'�
�%V��h�.�#����2���?M�7�Ȯ����=���/U�����4��2o.����v?RJֈG��
�=��%=�C^�&�R=��C�!��&<�X��?'����m���º�h�11��=�<6�����3�Z����@�,�)4g�!�͠�*��͌�ʯ�{Ŷ�|�n�<�����S_v��������]�P�5����%�Md�,�E(�]]mY��Y�� If`����?�͂ˆr亖i$����L�Wv�^69���� g	_yJ�=F��������*�$:�t}���p�/)K�5�{�C�C�$5gK�I��i�ܫ�/�t<Ĩ��E�g��]𣷅��Xp�u��:R5J�ۻ�g�X`��s���g�+e߮��9�Y��|�����t壙x̦��%�
B[jg뮐�y�����-}��4EA�xP��]����v���)��|��'�.�zJdS�+?#���"�>�����5H�{�Y#Ap~!�S����1�Yȼ�c�i<�\���9��nbzӽ�f�/HA	N�K�)�D.Cs������[�D��Fb�<��O|<bL�w�E;��Q�u�HԢp���2 �A9�pRֳ�ZK�L�.����9~��J��vet�f� ���(�~��:��,��-�"��e8	l�v�q��x���J�(hc��g@��'��x��"��[4�#����p�IP��ڎ�6�_�!-q�=��Z���{u�����0�ͷpGKQN�V@-��;�14T�*SjjL�X���¤�"�&�?����Tmf�@���%sͯL��$f��g���$�ֺ�s.��=�A��`T�Hwяm��S�1�%� �$2��2kȶC�b�D��	��\J�n�(�\��	/��R����SA%�Q���N����)|����\��׳��*���7$�i�Y�4��οD'�4��"�T���T��~m'���*�"KšA!���w�M�2�:�U���`k��L*D��dm��EQ���U��y@���n:���\��|�����,܇"�G(�5�������{�{�Widg�y	�Z�)@u�R���%Y�1=@��qH!u,�$�6A�B��≷�#3���?��j/�m8��M`zm`j�#��9��
����V���j�n�G��o���ܴ:�H$=Nu��<��#�f���r�ϔIʳ���&��i���PM��"��LVp�����m���W���ޱb�6a����ZF��@y-��zv�H���[X�q�<�ֶ��b��"�9����9r��¡����G�z�m)y�j�y:M̰�aud8 墩�q8�ݜ�?xk~��Ls����j�r|�?/C���@|�#�`�r4h�.�-<sp�ߋ��� 
��9Ԑp~�AG�yr4gg��6x"���1(��m�.
W�.6B�
��WZ��ДjT�&F��hg�in��d"UF�Q{+�$�h�8�H&�C.�Y�w�;�*F��͕�PZW��`�l�g�d��r��a1�{�S��tݜʴ6��=+��=�� )k�m�NY�E}^�^���
,X|}�_��Ippm4��F2	�eÝ(��'��l���c��ap9C>�ʠ6�� �&r�jt�m���g�u1�֩S� ���ޔ��Qd��ܧ�
̡h����K��ڈ,��F��3!��n�'�u[�^T.ɝȫ0�C�W�Z��/�E���^�}8ad��pnY����W��pW�ĸ�_�a�m7���)~�{ 8�ƣ����2@l�@,-@^�a���*P�
�*��::D��tO��7�`���kh�A�M���G
�F!O*�+��:A\�5: ����j;]�13��~��K�Q�Nr�|P��֏�����N��#�4y&������!�'�g�F�=�H���`��{�m
�,}PM��'�w)����"�'6F�d�����\�>�dE~�.�YvFsOU�ʍ8fuv1��K&p]��񖹸� W�7�~��S�^\.ӞR�=+If���/Yߥ�.?�[ \X�eQ��W3REAk�nv-M�,D9����Y��_��@���ɔ��0�e�G�ca�4zO��	�;�����Z[�m1w�6p��>N��"�2SX�o�.N�	�\���d�n�{N��Ƀ����Y����!�:��#V\���}+7������M�jÄAGbN�
��D���+U9��N�r��rEVJ_Kz�/agO}��,75�a��A{Un|ϸ�֬��5���Z� [<kN��E������j���׳���  g>\LJ�H	;�hΎ-�������*Q�\���� ޅe���h��"�	ܰ�҂*Lw�`%��-2vA��o�;d�Z���[���F�r<�?�&sb�2@^�����@�&�`���=�����XoB�M��986^�\)��֢a�{ɴ;RS-�bZ�]qg]�E����GH��v��(���Oa4?��P��/r���������a8�~Wf��^���l��D�	�9�8��������JL�HP�bQ׺<Ͻ���{~�og}3���C9�Ĉ���w��>�����z����ݒ-S C	gB�(������p�<�i9���2��Ob�m����WUY�D�'�e\��Jbm�i��j�@�����|M��ѓ��zWc���^R��^l���p��m5�m����	�Q�+h]���x�Cb�����F���K�U�����@��
 /��F����x�p��I��S�}K��a��P}B12�"V'��p]�ߎy)5�F�4�j���B��Y?��b�q�I�? I��Gj� hz�s�8�}m%J@�	e�!���F�:�� C��ee���_�^ܝ��Y��Zb�t,�����q� �W��>��2� "^/��?;�i�k����,�n �7��q
�,r͵:���R�,���]u f&Y[�� ���5���{6l�$�1 \:�t������8݅��]8<��n�`K>��E�*�	53�㿺��o�5�,�b
��z��|�ȱG n�a�S�]Jՙ4���I�(a[�<Z�VWԽ�%�kw��R�`+i�{��w�l6����}<=Y�Oo;�D��,�S� |"k���M��(0~�J�}����L�G)NC���A��ڵ`�N,�d�D-b��	5Bb�m\<��K�!:�VH&���emZ6�| �F���}e+���I��n��;��~�xϘN�Z��Y�>����q�4�[�h`؃-QV��q9��}7Zp-�.�a�C��?x�E�$}����=����:���4!�1�Z�(��� �qG^�3�7����i�#�ێ�)���k*����q�h��^A��@�^�Er�>ޒ�wG�����8d�񀣪�F�����FŴ���+Rk��`0�Ǜ�bZI�ģ�L����r�j�7��Ė�L��3�-ݓJ6��YFf�G:��׶Q�w���'���"��!��U�P61�>�`3�Kc�N+�ߚ9ƊȔ$��2�v�����,��o̤�ёS+�\���A��v�����0'� �|��������1 
r%��"ӦM(��(���^��.���T��	)�4�lw
0$<FĢ�����=�]��X��0��X'�z�c��K��b~u�9�}eo�N���x0���|8~���tK7\6�'<jR�y��H�33@8%17�X@��B|h��S,��N}�&?���PGq���ʫ�4w�g2K�M��Ro����ƒz9�wM���u>�ѻ����Cz�Z��8Dۅ�L@��5�N6R���� ��o\g�,�O��9G��y6�U�5�W���7�LOn��e�Ue��*�����sR���颾��ө�,�kXyq�_Z�f1�W���k��b�� �>1�8�DG\�VJk�(כ;��`�}�؍q��ς��PĨ�+y8}�[A�����y�&��BM!Uy�i��ph�pr���yNS��'Tf�����9��??�sȼ9�p�9Q�S�Y��e٪+�0���~4nc�i0j]�5�����1�&=�6��@�xa�S�nԖ<.��S)ac,2́"�X���a���V�%	 �Q��1�~*��C�G�yR�U�z���"��{% P�V$��s���k��[(�U{v�B�U��n���)qI!���jVr���������co�>h��//��p0V�h�T�V�I/^%%/��멏5�0�9?���1�^;��u���O|`�����`4�Ô�-GVNT4C��Ԝ1�'�ϧ墋���,\N�yi�s_��'%�d��v�N�,��nm�X��҈=խ�Z�����2���r*f2w+��I�f����1E��5�������4@���Y&,�~�֛}�ԽO�T�.Wl��&r���"����*���!ݧ�L��]j��-�1�U ��o��v�=4�6u�&,����e62��~K�+��*�
/ؠ=�4���_֨4�f/d&���p��5LO�.~�2S������Z ^xyʹ�%o�Krآs�Lj��x����\g�0�N�{y�KW�)��Y��`��nG_	�hgH��
�}�U�h���LXO��*��jj�˲�?�� 0H	�* �r�i�9�ǂ*O��k�J(�$ox�ug�{�$���Zk�� Z��B��X�Z�Rh�o ݴ97
'{Ir˽�l���������j� ������fA�\���J�����Y��h5F�w�_���$5�r͍��	�|\�mӮ��^��6H�]-[`�-?��]�U�$�'��G�-�@V�o�H�:I�����[��[)���a�d K�_��V��#���M�I��q-�[��I�����
��� y��#�������Bݥǖ����9}gF��`�\P/r�A�4���X6��ߨq�(��mA�Г[$
)E^n_��X��^ݻ2�wn�W�]H/m����R9m�M���J�M���}�#����á��C$�%NN�c��b3뷽�.�c��i�8iپ�ikQ�`��/�Lד�_�Z*�.���^t?C�'ྫF����-�yȹ��;o�0��\o���ânYGo8z���N��+6ɂ��,�x��BX�/�Nv����;8�Q����l�}pIwEE����X���u�N�.v`��Y?�Hf�����_t�R���=��қ�]�J5�L��"
���ٌ�MC<)=����;j����'Zg
�C��}3Õ�rxᄼ`6�^�hb�΍R��e�O�~��p����d�1�>M�M�E�<�P��e���Et��*�v����M��0%������f�gi�zrx/,kĥt�B�ǹ�F
�3�3�i|#�,��3�����͏�J���/���9h�ԙ=�	�9��ZcM�����a��/J^�Q��4I�epJ�2u:�a����AJ�*�v{�ߤ�k`au�/��$#����W��d���t�j�Xq�-�jy��<�թ��V}C���Cr7���cⶣl1�Z���M��V�v�'�ǛR���x����ژ������gS��x����/}��AA��$�[�;K��pi}v{A�7��3����ͷ-Rzՙ����1d`*62�G�?�Y(�x���}�����,w���p2t����9��� x�q�C�J<i���)�ݝOX�י�A��i�H^-b��&��8��n��X�d������<�MJڥ�6)4�Ո����s#*��u9;Y���`���w��J0�N�����8�w��B��cI����8������������flI!Jû��5�+�bb8�y��:�[I��l�4��?_	v�ڑX~�^�r�N�����'9���?do#`���M����ia�K�r.�%������ &��F�k��~�Ϳ|�ɠm3�ʽAs��:�d�ŎFO3�Z@��-z�mp#1T��I�_P)�EԻ�_aUn/(P
H)H�ko��g�X��K������Җ
v��%>��`=���/�`�R�MF@�G�����R�M�3^f ������	c��{ĩ:x-ꧤ�^7T�?�����ʕ�[H��B[��g6��q���}H[p����J� �r�\�����HK3�:��h�^GԒ�q,�����D�����D]��g�G
�
�9HN~~$v#{Y�Y_a;���<��W~���]��&3�5�	l}3{^C�2=�I��1��N~�s
H�2�A�<��"~�ᢈ
T�
�sI�&3�TGx���ӫ��;Zs�̱&�����������{��z�נ�+�y�W���ܖ%��99�6��Q.��������]�(�f~�r��'N�X�-�[�IN���8o����6@!6z���N�4a6�������c����b0.�0z��g�y�CDAs��ԁ��߻i������>��B��g/�����DR�j�[��,����[fV���$�ј�-���˱��پ8��t�W���Z�ҧ�ƪ��ۍ8TH���A� ]�t�%�x�Ē�A��Ԥ?��b��
���^��[N88�m�����s�����;s�tD�z���ܳ�����+�]�d�9�l�/xp�7\�ě��.E#FM�B�	~��&JN�:?�|�$q�eB��#�Kp���*�;�k�] �lڤѕQP��'� �	�����A��26ڑ��?���)5�E2p8%k�h�F����_	�8�8�0��Y`�K7� ��s�6�̞�I�}$��Ҥ�J���j��o��i�u�3�geO�au��o����7��<^F�%���"TQ���i��$���n���OЭ6H2���&�p�8u��$�#q��O�Z��~�^�*�mL� ���ݔh��s:�5:(�Џy�(����G��t�~�1A����<���u��Ӓ��n�(��q�!y8�&��)������j8��-i���5='�s��s�J�B�d�E�#n/��dg}]��c:{/�?xc x� ;�`)���^+�o��c�}��0�pW����.0������	4j�Q���h��L�^�Q��im(����P�/�E@������&�aq"Y��_��0��r��L[�+���s^Ɔ��2��5t{\��+[(��e��Q�f#b���[����D�Z`K�]�f��k�D!�n�b���l��iL�-�)?���R��3�#�� ��[ͦ����')ǜ�s�5<Mtc�K��4����U+���w�.�=���z�����p�}