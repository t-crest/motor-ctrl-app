��/  C���li����6`��Glwf�<�4�؂�˅ȃ�O��/̐7�C�g0d}�^�:� FkY��-#t�W���U#�e��E���$/���{�t5k![�4{�,��^��լ�7���%��~!H��_l,W@���3�%c=��H��f�%M����K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<�qן\DzS8o�렆e����rc|(����u��ϵ\������Ug����Y=�9K��:Q��H"߉���o����#�H��jD��2�@�@{�/+:ޘ�	-�>��������k�m���*�*	Ar���|\��*n�5Q%|��kT;�4�m�L�����i��m��Lz-@�����s��ƹ�Nr�Ӕ$��5���d���E*Y-�A5�r�h���!��C�;M��uN�T�jO*{�% �K���������M����F��:��R�����r)�ΰ�-����:6��@��c��.
{Fw�?E98���O&��9S�!��c迵ć���B�ك8?Z��W�^*ް��ʞ��-���H�~k�c~C�ӊr3���^���r����o���O�kPü2�y��;�������ȁ��+V������4�OdA�
�i��c���6E�1$�Ѱ%r��l����j�fG0>�
�@�{1�?�܎ӛB�g���i�����k}�㳌m�aJ�ç3>�'HL�V	C��ɇrN��l5�>ü�t��xW����*)�#��5��C�r59�a�V���}�����><��H�	���0��==8ݻ����Alע�k���:��zы�lɫj����R�49���"*{"r����|׃���dΏ�m�|Ȋ`�'�ޞ�cm!��AV��wנ} 3}/G,��wJ:�N?o����,Q�냪"@���e������>�G�� ҧܶ��K~��2�d�/��'�4~�-�u!aS���w(=ݓ,��L[Ey������Paо�I�����8W�m�oN���\��D�sʯ���K[jFf���&7Е��\��� ���}1��� z��E܁�UJ���-��p��-�^z�ޓ����taW�F���
�A�Y�%n��|��D�@�;g=o\��I�)�!���p�������<��T[	"��$����[����z?�2��$v�y����p}*uܶ\�x�pF����p�,��+�1nv�v�0�ڭb~���v�����Rg��6|�ؤm��򛁜_<����_�����od�����7�x	����,Opy9(��D	�ВPOU5��;��r��U��ξMO~��xO���I8ٖ�;���&��.�D�씩�A���k)yb�
FW��[�!G���J���[�I�e*����)%OgP3$Xv��(�r�J����I�xP��t�ٿ��87l=�A�b$����,�Z?��,z��WM���w�<Vܦ�kZ�MB:�}�L	-�5lw�w�i��z�s�>YZ�jҝ����}����8j�� �����:��;��@�N(Y�����|��a'�_�0��]O��E\%Ď���y�0�]�8��o����bc4�f}�F�_1���@O�I��^)��ԭ@t
Y�#{N�	nZ�y�Z�d�ڡ��ݳ�UU�4N.�C&���C-m`��@^��	]�f3Ĉ�h���9[����v�I�;�������-�a��EN���m#?1|C���D׍��	f�W�Q9:X����m)2��������>�9��w#
��`މk�'�i�4��m��g�5%�af	�ʃ����C�z��L*q��w`�,(�"B'0o��Җ�[VaT�S�f��ݛ铟?M.���F��=O.S���1}�՟}t.M ��������ė�8�ǐv�J�|�I�̍h�΅�*Չ�����}ǣX�#����p�b !8k�p� �����"Q\ے�'F{�	��.?{D�Ԍd�s�G:{V�*�9B�#�����s
�B��\YZbim�t���N��EI��>OH�������Ջsz�չ�S�9`T�<)7g��:!���|<sˍŷ�w�~e׈@9p�krͯ��<�6��󣠍��c�h{�����}"�I�&��V*�nvk
-�.\�A���� pr%���T��+��zOǹ��N��'$��l�y~��1:3,�'YL-ɳ<�P8N�"��^����iO�_��21r��<�2�H�L	�S�$�kRׅԪx��*_��v�-z�n���������� t ��u�Z��z0��±����#�9l�Y��9�����4=Ѹ�`|��I�x	��j¼m��������>���c� ���!�92�,�Mb]t����26KǢn6� [���Eon�6J�>��r���[_`�+N����,��������sy.�'��\\�㩱E z���H��T�+6�&;��W��x�J�����'I��E:�阘6��e�V7 ���W������9W�ښ�P�5*'«�@>�_��O�dKg㫏��Y��Bh>1
���̂���}�����Q�:~��!�t�T�;�}�5U��]��
t���C�k���@���я� ]�M��!3�]ykir�^K��"ͦ��na��wٰ<�ͮ?�ʋBG�ɣ0/Ѩ��'fe�$Zv��`,{"��i��ڬ}7�#ǖbɶ�����QfL�`P�<lXh��_g,��ߠY�7�J����)�(;wy����š�� ������,P��=3-$5��-��<ۄ/� ���I�rE<� ��0�� 	�	o#�'B�@В�kK��t:,7;�1нz���+�@[6�Q�������왁��K�K8��F��K��W��7c�W�Q��ݮ���w���m��Y������Tq߄� �gk���ZOX$W8Yl���kt�,�e�,�n���U'v��η�G6�ׂ� �r]:��$�)�M>���b�Z��x�o>d�t���wtM�jf�F��,��u��Y�k�b�#$������K�}v��-m`���*��6-��J���M`*�����;���Z\�xJ�^p��_'����r���ӻ+Qf�(J��f�ś�pc���^Z��_�jL��a��?M��2AY�7T����6b?�2�)�~��~ʶ�e�y���O806vv�I��d,
���u<��	�t�;�SD��|;��]5�C���:�����>s��f��^�eJ��p���U����$ʣ��NR�g��>�N�+��7�!�G� ��E芠2����#����y��PQ�R��G]rs���:�o�M��T 6��@�P���r��n|zF�h艺#�͞�SK�:uί
Xȥ��y�Z����}h#ߪ�~���n������r�#�+ۊ$��,��Ŕze��6 �����n�!��?��tl��`*�^�;v�3�D=��XA�s�������C�߆8O�%���B#���ҙ�</6���N�@�T�6Ԋ,�����D�{�OiE+�ш폘��W�*Z@̅Y߽t��-�s;�����3����}��W�l�}��,�Ae4�����(�K����˪���(������5�1#���XT.d�*f��'��2�3lcT�˕A~	�H:E{�3�a,]�=孠?��
< ٘\	e�Ȏ0
8�� C�����W{�U&�Gb�S�$ԫt t<��t�ѹ���>�Ӽ�d�z�ݎ	�y���d;��ƌS/Tp��	�!�vZ/��ʖ$��q4d���<0# j =q��-w���q!�{A�����',��N�יW��g,+�uy?k�+��a3͇%�F��kGG�*����5:��3�l>K�YyŬ���`W�0�-�+␊���^_�!��M�k���ɛP<�]�}�lԑ�	Z�p�PO'�����E���U;�9�ܟ��1	m�H����~��wh� c4"�lS~�S���)���
?�|i�ygw��a�^*��
�f��X��"��W}ܦ�9��C�`�|�Q��lAYhX����ܒ��R":g��MЛ��,A�N"!'n�m`���쫐Ws����7G
�Ŗ�C���@o %ȿ��95mH����[aY:����<[��m�2���u�3U�h`������?�<��