��/  f���1����o��%���[� ��w��^s^�����q�6c�BO�u� ��7p_�;aCS�㘕�k�S5�#���>�R����L��x���W������9���](!�TϿ��Y�
��
���B�J��T^*\e�l��<�/<Y���~�tlz�O9��5�^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK ��X�ش�[\��i-n�I���G��N��+\^�� y�p��PKA�!�H���kI��	&S�I]����BR��cs����&��厰]|��������s������wD�mݯ�?���ёs,iZ~1�=��z�.��oۓ�"��a�p���}>���MWVF�!�a��^��i+gn��fP����>�{��T踙��r������U�����E�H��(f9��.ϬS98_���J�M<vN�4y��	��4�#O6�0�s���fCXBA���4�z�ʴN/v�|���π
���O������T�ϯaxU����S��W]_D��E�1.�TgZ�h
	u͋�W�Xݜ~��_UP���8wg0�K�rA���_3qk��*�>{�&؇9��'4���Oso�m�m�)��hЦ��T�m��e�:'(�c�n�cE�8��p�f���3_2��R�2�"QlV�k�i��hN�NU��t>kKΗ��9?`�jK`�!��Y�#r�g�b�մ?��>���.o�t������M�ۥw�D��s����^m4����i����w��/��Q[�A\\��� ��Č��/ 0��(�tno1��M��xi�V��e�O�ǎK�_�Hgtq�J9ҶO���6ɬ���ٵ.����K.9,[�[̚����mY���Xu�B0���P+j��2��O�Ab8h��'�]�t�21F��� �8��@��D���ņ��5& �\ʣSTGѼ��a��N�A���:G#j��P?na���7T!bDFY�Y�� �&������ռ�Q0�/�!�E\�q� �����Y>w,�j�]X�0)�2�{$ 'ɶ-d�a�J��ŋx�RQ�?P_XvTüM��ڛ�R�����B?Dӹ�R�Xu�EGj���L�ULKm�6�������2K����E��N2��պ�	@�d/�ː> �cy#�2B��Ӽu��_�az�D���RTRP��n�!��EZ㦄e~�G�/qɬu��=J�[�Ie���$�Z.w�/���~�5��;F�k����b���j�b�9.�h2�ƨ�@���,��>��`;qŹ�5�8J����u����o]!�����a����I�`�a=�~޴���Qx�7��7��������E�嘠����n��ۗ���-ˎ�+�7sHd�NA�~FJ�^/����Į׃��2j��˒�n����?�;��G�J��A���,[�=^� ��u�d�9��Ҩ_���u�i��� �t��7��7i�=�?��9��ێ�ێT%��ǡ�E���kg�B�㸼�{__����?[�Z9��Am�f�>�h=�
P��%X7��ٖ#�s��=�*Su���Y��{L�m�Bi|y�B�w��c��]Ի���AV�wGw%�C������{����u7�U�Z}�zoH����伈b��×Ȉo(d���Uml��q�s�ș �m�`�`,�E�����U�3��9W�&����A�FT&㙐��|_��aa�'���R:@�K�<G����Qܘ:j����@{9�N����$�}5�!3 �1 Z@Q���X�����wnA�����Ð*����Ix�
Y`�'|e���{�LPw]F�=�M2���C�[���J4�z�^��aPS����H�B�5ZKG���5��K���ԡ��+�Hjq�]̺^�v���w��@��V�Ѝ�R��7@�LM֛,}�DٵE[��ȴ�W�+ĢDu�5A���m�������jm�d9�A����3�����z��·`���jS�&sr�Ó	8w�u����ߺ�ʈ{Fm<�Eg�y�����UIt��daCʯY��d��<�n���ЇM������<S�`Ʉ��VD��&y����d�W{�,7Fo�~��-3�����izRL��%�5ubD4���ox�kc���ˣ�t��ǟ�XC�{�v�~]'a�u��]pgg1���,>�.}r��>����΅�������3n$�\�x�%�,������{u��0�[�s��\���ѹ(�5*D;1�pm���30Nf#�����2Wʹ:���"��6���c9K��e�O�'���5�u���"?����te��L�G�@�n��m'5A�aO�{d��"/�@�c勺L�7{�+k����r���>tƙw� �n�
1j%9.���Eހ��vn�d�C¼��������k^M��Wk�P[DR�NgV)��lw��@8���}��Ϸ}dZ,�|]5Nv��sa��:y�/�f_���i�WDUS�N]����e��`�]����ԅ���j�f�
OPf�W�����r���-�§���i�|Vp����=-�PR�(�p�%e,�]�T�,^�}qX�pj����[����M�$q2��/�ɞ|�6�9na��*>��|9V��,pd%�4��@�� i"�'|D"C¼Aß����ס8����o�yQNp��^�9[S���
���*�T/@�iˑ�"���y�zC�Q
�lw�&L	�6���V0B���V6Y���䡏��m���v��q2�&̦�{��u�=��c�а`:����%;��pQ��,0E��B�� �m���}�=y��rRL���*�o/U8Ѭ����౼���-����+d,{d-�͵��fܟ�*�E�pG��g���$K��S�tz�}�,���3R#&?w��$ś�ğX���C��xj�-m���C2��'7�����K(��Xel[P��=�J�bvM�'[���``�!���ﱬ��p�s��rDl�칝,a�*��}X���5��.�j��{0+0//�^�)H����1���^e�R�`NIM{�����,�c	|��"�o��fչ�}����]���WJ�\3��=�c�tF���PS�Z��M^I�OV��#C�+��:w��o 5x���永<�!d����V
�؆�g��<�"�vb�Լ�p��7Rc\U���/O �\��
�X������DE�.�n�o�0B��у���fp1�ޕ�ᾪ՗ѭH0p_�PYIFi]@�^w ]�)d`�/��3WCp���
�;��untc�o����Pn�^h���k|��!:���E�MG�L?�wז����&w�l䟳���Ա������pB�]V���&Ux�o��_~dVl��;���<-��������f6�p
��f����>J_/��22躆�|�d�i��w	��?�E���� xM�+{N���ς����i�ӳ��0���B2\&vm�����l�f�i�_I�r"B�����]�x�w#@SmՇu�s|�\�IBp:~�&��o���}�Q��K�����3����H��ƹ�9D��ȝ겡'3D]O��aZ,cq�8�96��p��٦��M�����(�B�3����:�V&�]I���XM IO6Ϟ�&̸Y9 !Ҽ^�K��Z��BUA=*��|�K�O+�Q�%hpL�d�9I7����{V�-�T��> X/c4bЎ�S�2x�����ȤqI�~Y�
I<�"�L�蠜��7\G��~�,]�E�ap��LX cUmM�8���jBW�Xc��|ݬ"h�$�/D��e;#���gjp&x9�����Ұ�|�`oJ��;�,<���%:N �-�qn�n}8>�5u�w8�3���ʚUﲖB�������ҤZ���
��g���z� uj��� ��5wX怷��U)C*	���*�6dܢ���g�͘�xm��tT�}�h?�:@'�#�	{�L�))���s[ɸv��R��lʊ��xeJ]�`U!���SyR��>�O�W�8���+T���i8�x `�[ =!�l�����Ü�-��O�����
��nB�OFGK����鲀 ��!ra���f-1Í�"K���l����y]���)�v<�HT�c�"�* V���I/i�2�xgB���	 ˋ@6����k���V��	����a����<7?�^n$�۾.W�@�w��1'n?�ϧY���&�|�5>�
>y�+:�>M[3V2�q���l��
u���$���� ==�k��,Z��H�*�Қ�AH��p[|�k�۰�0m]QlS_�L�����A��]��vj���W<������	�U���Z�ǳwo��8��
�ć�Ց�[d��QM!���!�K�7����t	FK��m��i%	uc8���Nfd�����lo�ZW �7ӂ_����OҤ�7ۿi��=D��������/)�x�6{�ow��n��KD�b������؏ PFz;_t�"�6�ܰSC���AF}kۣqK��S�%ƖY�+��n�B�f�ƅʞ���h'�4��̐���Zy�տ����9�n׾Z��]��Ur�RN��տJ�ܽ�]s(cP��TZ����)������J�#�{�t�IU��[2(�����mv�[P<�<F����w�P^�	�kS ���\*"��Y�Үdl$������2ǚ<S�cw��7j�g}A��vֿ1ٱ����}O ���ߐ�q����	����+($����g�SQwP,�F\K`�
)_���ۅKI��HÓ���$Hnh�fw���*�O4�=*<���VΞq%K��QNY�����5l�D�&���{QY�L��3���^w�~���@���$,��Jl �k�� y��IW`���0K|�����-i1��Ji[����Xq���'WȖ�����n�tZ���C>��6]�|���̼?A<������4�w�(m�!P�BGw��S&�Ѵ�6��^��,M�]\����p���q�T�O�y]���	6��V�V�Չ�5�^�.�o��ߜ���c�_^fQ��K��N�5��O�yU�Ç��3Y��a������M�;��>��}��cT�Ljd[��W��
?E��q�NV���v'�v�����5�7�������}C��ոK�@l�$��b�ݖ~/Ce����V�¦*�\���k� t�S����ء�?g�X�{�颌�MA�<x������'��s�)}`}�V��r�A!1�#b��D�m�֜R���U��+�͗�uz' �'&io͓"Xܳ����0{>��z�Ҟ���V�#bC�Q��b�N&��<H!�!���5�h���0��%���W){3y��>��r��ܩ�f�R������O���y ;U�0�4x��"�I����f:ϧ�c^�AFu6���闯r '���t��E�9�B����=J�	��:]�3�n	u�[�9?��2MY��4
�C��X�7` Q��
��e�7�U��5��lGT������H~,,u� �R��MgC�����^(m��`s� \�'ر�_9�O�	!�b)x��Yw�]rn��Կ��n�{�򖨰��e�c��9Ŀ���T��;IXFT������4�,j>]�E|焋�}�@������f��ì�!mG�����NM�k�@2`7��a��5tqQ._���+�}��>��A:r/I�
�B��pd���t�q��"v~�W����yF����;�4�f%D�E��g��~�{���0|Z��	8��S���9xp"y~���̿�n!R�y��
\C��ٙ�q'_��*ǟ�RЅa�$h@���ј�p%#6))d�1�58X[���#�	�+X%rX��Ly���~�]T"n��{����`ৢ;��q�u����Dj��k�����y:߀m��pI�84�(ZD;E܂xKOa���w��W	��1�����%�Z,������]y&��b�C]M/:����F�mnwE=7���[�S�y3�/�yZ'�Č�I��_`�;W��J�Z�������2������)W��'����BJ��G4��cƚ7�����[��+��.�	�FGm5ׇ9H��W�l��w۶�c�	h�+��|Ѥ�ԅz��I3u��ָ���v�������$hy@G�O�ֻ�Z�r��FJ���้�,"�Q%.����c*B~���9	�c�B�D