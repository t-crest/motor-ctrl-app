��/  h$�p�̦k�m�ٛL��?�t�N\6
PX=r2 UV5��jݴ�vJEB۱��#�y���6c���bo�gƗ��GF�N��Xʣ�\L�a^��8ە��5"��8��{H��\^o�L.@��8����L����:^8s���c�{br�䨑��M��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<p�at*:�I}T��3H����mi��$�+SVj7:�����֝��/��%5��S0Da�I�`6�?�+�*��q��p|�ħ7P�9���8�Ҧ3Ib��i��F���3{pX����
q�A���`ёC��%�K�*	P���x��Z�7�T=J�E`�����u�ֱV�K��T��Q7�j�SQ��r�ٶ�ɡ���ؐZ	FN<���o�3�YCŏ���lVެPA)�����C��0{�sZ��Ԍ)�'ʻuNO�o�(P���6'՞O�l�P�� �]���I����K��?њz�0���zTPcK���+Α��ҍ��iB >�z/�"XQ���M�4�[�#�\�onB���Z>�^p�y����-�vGrE��a�/E�)̺
��&�)YGL��Q$��Y��(�D�Ӂ�E¨��}�>�$�aǶi��PO�Sbv�o#h��x
�����4��f����t��E�թ���L̷H�������Z|��͹��I�d}Ѥj���*���.p�Z�6(^��-��.�+D�0�� ��j/C���{�M� ��\�O�I��Osw��8��\�5�&�D3B\i+k��"�|�;'���;]�t	��b	��j�h{օ���S젡5�,��J�6͙Ӡ:�3��ptvV��8^Al�R�I,
Y4E�b�]����j�i�L��`;"�}��/CafTz�ϤP��M�a7v���] ���mjhɪl����7�*�~�]B������!����ys:�ʌ$�f(v�������v��¡3�3��x�ֺ�kd8T$��V�*5�M���R�~��~��Wc�>o?m�@"ӓ�Hٜ7������CnU�p��+o���)�< q8n�m���8�{��:�<5���i� R��\�ܮ�<��	
c��G�(fC1ˆ2X 26&/T����:�&|�k�t=��^���Ě�'�.P��/�hB^&S�&Q�M����`,��~��̎�u�5Tv�x�=�0/�Q���>4F_��b+���v����Q3���ػ��X|�������7F�r�z�Iki7��s۰G�m�����~�p��z2ؠ3��iy�[�8ڤ�D�m�/¶�]�Mq`�K
�T��_�3��֧'�d5��)3��j���i4�"�0ڱ݊�wr�����<�rUF�9��D�^̻�S&����?u䎒��.%Α<���2 [.�4�������&�<���漸��t|��I�n��J�P'�BLѬ�ڮы�,��tK��ʂ�)p��,wsqm�|
��p3'ݡ	��� �O�`�^!W�2�J��84��ʘ�f��F�e���(J�d�Ƒw4�EhsZ�Q�
��x��Х�_X�Z3�����/�?HO��t��$�s���V�/���x�1c��@��
k$	GQ���m>\���`����#���Nwo��J=mb8y�(�;�#7AG��8�ď��1�n:AϽ���X4J�]Y.YC�g�)�sO �4�O�D�>�dϳt2[l��B7�G�f����p���D�^M��$��?;�������Ks�pvL�t���2me�
��E��#{�+¬4<̿�ޞ@�>7o�Z�E�M-2P���D
v��n8�Y����SG���"�̀�T��y����� U��r���2E�W�O͕D����Cr�WP`��'ק5�~��rT�'�[�wgm�]y�nE� 7m��M����ȋ�9\~ewAH�ĶNY(��pvS7�|�Cw �m1�yD��;�4Őd�������%�DP5�2/������������H!���uA���2�W��(�PnY�h��w�E�<�`D�0
�cm~f�w"�O.bi�5�ԕ6�jAMwk�_�c���k��Jrעy2��:|7���r��Emu��!���yʷS`]�� 	82�.4����,���"M~��;��������{1�Ic��J���pX�/���1�a>���`P�/�����r����@��']�r���E�ñu]�%���Mv��!�*����q�1�BJ�p�����w�+; �ĭ�)��	�h��LZf:I��/�:�UpM��NlI�J���)���%J�(j~��gL���H�Iy>��N���Tc%ɻ�v\m����n�wyL��'���S���u��?��zk�~�� *"��yp��y'.~p�fY���'�HF�����f2em��n��=��)�s�3RO��f�$,x�V#������ݐ��{m>�}�B��|=�U_s�1$Lèh����i���u̓0�'��|n_���^Q�$�A��num��:���
�J�:��W���}�n��M���٦�=�7}�ª\�߻L*�����g�ZX����R�+��E�;�|��Ӷ�UH��^]F��>��Z��+�e�W�T&̅�p�i!�͒�,�/���a���X��l٦��{�v��{��Y�X��� '�HJ��D�CA�'8+��@���Q0+��v� ��jU�)&Z�\;����y��C���]#h[��k���-�V���<pH�[@u���{-�(��ާ-a'/��(��:vт�E�r���;wվ�Oj?������������P	�0us���ĳ�4��-��A3̌:�&4����q��je�>o��at7R4ќ-+����r�?'�9*��ap[*,:���(c����$BF�9{�:Wa�,��1�@�q�b+����ړ0e�=\�W����x�:Յ{�(8�oڠh#Γ�%���� X���"&���>"þ6-�=�̥p�����4V���ωO�y�0 �g8��\S�w���|�Z=ˉ���2ʠ���L�І(����ĸQd�Et3�_������e�z�8ݔ�t;��֟#���
��B����ȼ�A�?�r�:FF�V)B�H�Y̒J��J^t$v��%BI�۱a�b�vq��#����_���j�SC��U�L��kiעSo��i��bT�#`���g��yJ�PaP��"��MSZ���&1Q��&�������\̟��o�����J��>睓�0�؇k���MQ���y~Ͻ'�0���&�b�*Z�=Ef:�qW��?��Nq�50�|W��[d�p�Ⱥ���eU�Ha������8�O��x�9t �����}�O0#.&�6�rW�����>���y4��Ք�����gz�>M�:)�KzʆA�C�2��?Ϟn�<�N�~��Y���kj�\����|�웽��%Tfh�GY,���ש|ؾ=��p?�n���b�����>�u�*h�(&��m'���A���Ѱ5y"N�!"Ke�{;G�K��X����P3��t5]`Z
d�1���Νɧ!	�Uv���V�&z6Q��I:�$�il���u�j�����{�=��ޱf,܂�p�#��y�J��K�J�PP�f0v<�t?L>/	.P���8!~�,�C�0�Ҕ韟�2Bku@�m�H0}�F��V��ۣ֓��,Vp�&�FcgI���Bf���04�5��&�l��f���d�Nm�Z�j�s͟�ftis��O��7�Ά��G ͥS�̷�$ɮ��ss~ݩLT�ѥ����uQ8.�ܝ�%!�F��98��*��������� �*H�}=Rf�L�mQ(��	�T`�:�Ԃ/t+�Ҋ��D�z4c���VY^���̸R���
�v��5��.}j�f�w��`nF��}<&�ibː��َit����J����/F���9����U�ƥ���]�3��o�:�Dt��|�^���r����i���ͪ��	p�vl#=�/��8b`~w�{ >�_M���#��jf&ɨ̚�<���������¯2K�uaa�����mv���'�|D�O�V���?4M_k��p��+��A�֫Wkc-9����9u�V�oPQ
�K�EbZ�a̩�4�v��z��	�������3!ԑc�S��N&�1 I-.v���)����FSb��k6����]GxAs�{�9��'���˲G[��o����X~̠�y����� =��',T�5YJ�L�[�/M�1D�Ďk#��:���cs'��{u���\?��H�q�hB�gJ��7���U�W��oN��*����c�{�wT�ѲB	f}a�Q�=^��� ���ĳ�0�����bkg�W\*5w���9�����*�- �K�X�wt�V؍oT�D"�{�Ƌ�c�O3�c�S�eˤ�[&�̒z�X����D�n��"�q+,�ԯ�)M�d���'N{)б�qpf+n�>l����{$M5)��e�6pޒ���ٷ*F�f�A���"��g ��%�p�.#��AX��ڶx%0�F%���0u�7�bl|�EV�ּ�H��K�l8��~��J^i���
]\)�K��9���C#Ԣr�`�H4fq�V���%�"ٗ���T#���B�Wp����f?���/��.�����g�>�To�(s�s�~@�[)�3�51��8�1S�ב7��N���VZ]� ���NMW?n��~��p�X'�'0��Xe�!+Y�}%�Z���/*H�A��(&�
�|f}�)��y��|�WS��5����GY�P:|�x!C�GU\���֋�w�����O�7�&�~�U��<,;+�Z����dw���5��6�(ԩ(nў(���Ex�5?�Rp��K��|Z ��u��}���Aq����D�Z ɐsR�v~Z�ڡ�S��@X���o���H�Z��}m�ǧ��G<v�󿁽��RbR�|��lc%��c[�2��q�T�lG���6�cPLl�W�y�%�dL�����s��)��*5Ԋ3*�W���i ���~�pa��7+9��yh�}S+�G<_)��
���RLUgG�������
�fH�����ǿ����]|��	��~v8�si��3��T���N�x0�h���_�S���h�8Q��j�y�@�?a�V}�W�~��q*��DR����Tl��3D2�[�,����Iq���2�-���)��+���ˀ��*mXx��@����!ͦ�L���m�J�i�>|��C�9���9���	bY��Hc�Ob�)
!#���%"Se~ؤ�2�	���.lK�g?�*/~;�P�3�-��<�; �9,��V�X�����e��G��'�01Q��*	R&A�_AFP��+'�5��c��r��v�*E�hy� ��͘>��AD� �d�z��*]@�!��W���f&��i���Z�J;�ѱ[��?6�=�ߣ�<�-�Y7t��Scv�!�1�tG�� ,�O~F�Vϕ���҆�$.�w�f��<u �]�M� ���m�pu�������7��Y	
2nG���ݠf�eb���`�1�,*�OM�y؁0�>��=��I�]��C�]��]a��<r4i�pCF!�߿z��L?Y�U2D#��2`z�����:yv���yO~ɚw)���+������%�ת/_L�s/�w�P{� �O�>5�V�!ͬ1�pDN���+o�i��Rdb����E��)xQG�C��9ǖ�08���%�'Ywq&���.FCz�X����A�u���r�7�Fo�_@��%@I�*~����M����Z�o���n���i���l���-;�}�J��Aw]�T"#�f*>�G�5eD������FB�Dm1�ʄK�ҭ�c�;��E�i/̑&�2�E��1|�_q�Ai�;{�p�c/s�u�e��<� 卩}sm���OblK�H��A����XE�~���P����hSÎ��\w:�<4�M�=+��Q�� SQ����V�/�|+�)5��?�����E�-ZAq�wj@IU�4�	h�$�7��R2oQĘ�?b���D���Zz��.����,%�.2�Ts-زb�b�#�g[}�-�!����b� �4Jx� �N_�6	YLj%����$�:�ƺ����+���RX'h�H�� v��͘�yi	�0��;/Y���J�K4� �_�Y����U3��?N��dT�󾺦z���*S�QN[]6}:O��6�V�IT'&��'�g!{E�b���Es���H	�$����[�q�C��^@�$i/^�G$���j�n�*��{�a�pCt~�,AӇy������ߎ����jr��<���.��8��N*�	�0��{��`�w]o���>tv��K<=�Sx�t��ƪ�YGC����30��"]���XG���5GվQ�o�P�;L"H�G�B�j$M�̍se�(�v�7�K�(Ё�_of/���@'�Դ@��C�!7�j8Ɗ�n�w�ײt���s�E�l���(�Vo,ع0�r�g��;�<���&�'��G1�a(��Ԛ�Rو�}���&�|��SFaO� �o"	���Z_iDI{�#�ɷӪS�1�ɘ�hČr��+�HЫ.���t��:����`ZR쟴�|��y1j�zj�~�.>
��\�旧H�RQ@�ubh��F�j���2'�	J��E:"M:��rn�n�ru�~��AoT�ս얯r�]�N�
���*�U����K_
s��@�h�)ru��	��8=E���_�����7�m��?T�\�$���/�L�o8�����j7w��dg�*�Q�01�=}�ۡxO�N3�UY<�S����ļ47��q�z0����/����K���T6�B���Ki�����w����_zm>Ə'jt�BcWMDaK��{�T�&�e�8I]�Զ����N���^yxB/��~�`�����4M����>���0� ;�ӜʞTd���y�g�G[�R,8B'�E��v���tP�VS�,?�5�j�z��E��H����L:���ꎙz�V��>
B`Z0╔�����֔J�_ʗC����c#��>*��(qG���9�Kx���ȫ�]��J^z���Nx�%��%�?,��lY,����w2�ד��
ǉ�3Z)�`��]�������\��B�z�C^W03�Wq��x�8��h�F5t��H�=L�z����6���ܹ������%�f_�������1��fy�P�����;�CB3�t���]��<�[Pi�?���sm� f�{jy"��;�Wz�����O�$��$���Q۽#!�}� ��yu���%}T&�	E.��K� y���>+�ۑ���I|�\��T���v"�`J��O%�췡�s�a�+�Rď����A�S�D\Rʚe�*��/Ee��q ��L���]�T�3��=6A}�|��W	��"��	¢����7H��+:ɡ׾�[i6�krC��U+ ����f,~��q��O5����c�4f�o=�G���0�v�lm����v��A8��J-J�s1'�<�5���fD2k�q�h11�Rٱ=�����ޚ�>$���|s��n�J��X����` ��*�)M���c�/���j�]��&K'o+}2������!W���Ѥ�T7Ƙ�56�#�)��W(`�+Pm�>��$]Y�M�s�=B-���B��5��l���(����z�-^`'":tӱWӤj�Ǖ�c��4����4̬�c��&��~*�_Ǥ��	�`W�P�¢ v�>J�\o�ɊȻ�����TH�?>Ord�QߐԵ-S���*O}�5T�&mC_����W�^@�{��Tb�<,8��(�L\.S�0V�|��.�D_^S��Cǈ�l'ωƍ�����_&�uMs�Q�G����� <WV��lbw0�#�`�L�����if��/K���_��kq���[�/�Rx�D%�g2���'���#U�"�[sNiX�8�F- obO�8�^�}��Wʿr��r�?�9���m�F�	N���_Lr� �����������4h�wqK!s��Lc���X!��z�O��PԱ�m��
��R���i~���b�?�yXr7,�?�n��m��5��;\�%#��5Q�y��V�O#E���
>Ζ���{S�������PgL���0���b^�8��J��:yb=�r�Df݉����</e����}�f�9�\�wd3DH�dp.���q	6��%����`���e��G�'���샽�O�$](5�%቎��F�f�����Q"_��/gUG^�����g$�>�X
u�߼Z_T���{��[��rڠŸ��.D�5����8��I�볳b(0�E���_���¥�;Z�p
�lo�[9���f��& �DF��t>o�>���e��{d�:`�d�x�Ւ�����aH�%�eaZ��@G	Z��:c8v�j�m�:
-���}=�_��"���#��L�&�i�����!���6�3�'fh�O)��7��K0qr�>�P�o�r�{�k��R����%�ؾ�\�%&�,�����?�?_��l/�����u'��%��?�8LX�v��d5[�Uz�i�6���$)�Y���B>�~1N�ʞ�0R6����q�W&sUQ�Y����$�z�PE���AT�߄�-*i5-pu�`�w�Nk��Q8$�����U��{�0�^��!Z4}��������DH"}���p0����HS�F;TW�,��H��0�'��^ �r_��:�ZD��wpp�"�����;�����X�ܡ��}��-a�����ld�`w�_WY�Qk��+�o>��JƔ���*c�b`�4��2|O�Q��]RvF�1x��G�P��]�j�= 3d���S�C��l�����Oс�=����JB9a��3���Q*2H�Jo��Ϙ�\t��@��]�������|�b��(k����[ �؂�*�.�Z\�?��6A����N~�^������5����5HH�?��|��ǝ{�.���� ���ۨ����d�ț�>�E���w����emNR���t}�lF�L=n������A\E��7-�A����6�jp�Յu�0hg��>f����Ӷ�]	����з�o��}�t2ͩ-Xl����의���h�M~�g���N��1Cg�>&R���Q����WѰ�	2hn�v(�3oLdɔ��[�gEQǹ��j,�Mb)ʚ��T�o���ێ��aH~4�N֏<���?ѓ�M��[�D;�^�6���o�_;gUM��'�>h�rc&�f�����`����r.m�Ϲ�T�+�f������u�p�Mix�1��Y�v���֐�8Qt�I�atb�A�Z�$����`�`2��k�o�}��j����;�F���S2�4e謞r����D�N�:TFz����:��1����'Cd��
�f��V(@eY����5w B�� �I��|�F��%�l̆�UQ�����y�Da�ei���c5�)E��%s\��`0�����_�����VDxR�J�W�',�Y���N�۵���s�������U
�OƬyH�sD��.��q/���K���@���;G�*b������L&��n��mZ񏨱��gx[����t�m�]��X��� �y�
$�h\i>�#�Qݫ��?0��{4�~O�(�)�ѓILkW>˞Or��sY9�M����*[���f�/�D�T�[��{8��;:��D�6��=Mu�c�([�5"x�?gB�z~={�7�6��D쾸7�*J�|#��V���I;��T!�pp㓥~��i�<r�6'��F�{��E�Fj���*��uz�*6*���'�����[����������z�W[�_�ӫE�?P�d��[�� ?3��Ԝ�"=��L��m}m�M�#X	!K�o=�>���c���'�C�>��boL(��Ϝ������ۑ�5�Bjm<KOZ޽�Fd/�Y�Wvѓ��w�t���l���KR8T�+�ǟ��M�މAy96Ffo�|���3_�#~$M�$ח	�B��_$>l��@z����Q�`��=�sK�M�Q�rD��ё��=�&�M��=��<�X9M� v�ͥ�� 9��ԧ�N�e؁��5+*٥9�����N �(X�G�Du�r��J�Gr����6.<�e�@�r# yc�w DV�����Vi.�����y7����?2�K��M�M�'?��T�H�M>(6Β�$���NJ��8��`�Uq �d�?���򪄈�7%a�_��lo[ذts�;ץӖ<�JB\���:�\�=��Qٵ�F Ҥ^S�Z��Z�� ��ʧn���3�9�?�w��p ������	���'���F��V�?�A�gO����B��[ul�������7�]fx���M�6
7^�������S^��mOo���t�m��c�&oI�)��VCf�%��+(��S��X����q��A��7_�Z������KM19�
�<���֣Pf0z�ʬ��τ����I�K�\��J�q���OժQ��u?����ꏟxpgW{��Ke���%`�6]g��a[+�U4�?�����ɕa4	9dq�	W�0K�窧�YYD��K��F&j*�aq��7F�|�N��������,�jpO�u�����e"J(/䴞k#O���
){B*�4����h/�wl@
�S�0 ��׀�AƤ��N�ɏ�ȯ9��9ss
Ǉpd�)]�b���|����l��%Bp��%�6��`��
hݒ�e���⻖�.�N�W�8�d`<܂���"���:IIp��y���󍨗� �}OE3�ߵ�K�Ύ�
��y����y4��ΦI�)��QA�[Z���v��;IZ�+e��̍�yX��� ���J��N���g���o�Hު�)fV�����ٝ:�Hk�D��ژN]E��
����l�	��}5,���=�,?��E<"b�c�R������"����A���H�0}ȕ*mj(>����r���Kl@L��A��Y�ׂ��r�w���G��w�m�Q��nCbl�3R�+w�u�O~�>����|�(�t�1(A�r��u����M�A�:aQ{�˅�?�0��f����XLt��@��A;<�̞R|jŏ�/��;�d��q�Ӻع'M�_d�SN(�tX�*d;0X��e�º����L��g�3�ikZTs�wF[A��wK�$��y�z�����_�O1�j�Lv�t�gQ�V'"u��M3vm�C���ؑ�/��� ����c3��f��	Վ��|W8B�:�n�PT47*���^-��X�`���>�-��/³!k���CT��F��a��#Z��\^����U@,Sw�?��1�H?�֣�;�2�e���-E%	�5�
g��A�sj��1���������:�_�(�,_f[h�{ƒ'���p��0V�9��&�ΈyoW8K°<3i%�)��U���꿖(�r�{��!� ��sN6��<���IE>����gX�.�v��ǃ�U��/�BuId��I�]�6WM�Ǝ�~B��o頎a�`��W��K��R49����������.#��ӯ�4kQ�׼�>�V�=�u*�p�����_uKM��i{x�ymտ�rQ�A�}�W�}q�>�r}�mn`刖�̊k�&dkI��1Ė���S}��k�w>��I�l�	Ƣ@�p^�J2�@V����ؖ�$5Gq?�e76R��PfuB#'Ėe��x]��J�Y8$N��� �l��>� �/�_����
�3��e�u�ΐ]��-U���Q0�gtZ9
�y�B*�,} �g/#��y�bN��6�c����{���՛6��YX��Z_��2�,��93�HN
VV[��α;l��pd!���D����`�ը��kIE��D�����^%?�O�ҝ�g��ٻ�S��3��Z���xA���Ή%�v3+i�l4���ݪ�1�A��Ϧ���D Y�A �|��f�8���g*	�d�u������ԙgS�LD�[����l_ya�i
J���<9���Y3�T@\�������˖I�������b�I��W����%Rg`'��"fFn��?��u�p`��9�����CR�!�`Vᵦ�VY^�봛1��S@�'a2m�ɡ��<�"�"ô�E�ԻY���w��;��i�Ԣ�x���ls�0���f�t.%-� �YF/�Q�
 E�N�4��U�p����l�'GWԢX��a�R榳�8��>��b������D��H���Ӟu�2�/C�W��Ñ_�̍(.����(�b�PQ�҆#^�SǽOo���*�ekWu�	�;Sa?;��Y��&Da^(�x�K�{庑�8�M����%���24�Z$�r��ۺ_A����6����vH8SM�?��>�&Q�a�3	�I�
��L0َ. �z���!q��o��hQ^kuz�8z���+���)x\D�ro�k ; �й+5
4֖M���1�,�Z�v�G�ӣ1o�mt� N�^EW��C��fv�"��IG�|N�<O?�{�����XL$Dr�5`		"w�N<�Ex���6�_;�n�����3��W�;��.���0N���x�Q��OA}5G�"G��x`C� �p�<KkZ�m|	��	�:I٤�l�ʣ	f��M�R��kWqΕU�W�5������{[zjW�~1P�4�\����f,�B�n������Z�Zl�>qS&'���'��e�4��3 �9i�r���o�_���qZ��iɔ
�P=^�$x�������Hv+��(�(x�����nK���4�׻l���<(��}Բs,1��m�C^��Fd_e
�ʔXd��^7���O(7?I�o���ٴ	�+
NQ#�'��J��oZ'q�
��[����Ѫ��XI�
X��������.�@3��p���3�q��/��N��`!�
���4p��G_��I��>C$ߍ�*�_5�:={*貎�`"�aa]5�DJ�R(�tW�ҙ9>!�|���ōP(.��3����4��;�r����8��1(( )4���wǯ,��e|c�����R�M����#ؤ�#='�t���Ϩk����6Y��Q̊S,���{.b��ge�A�.!�A˻߄��]Y�󇦛&(Ǌ�g�>��k8�b�د�dv�wy��k�u��a3DIw�>���G��v����W�fp6V��´��&�S�,�@�qo��E{�٤�k~
�8�3��[�̌�F�0��5�Dd��D�i<�������KP0�_F_�h.�>�*M�S�|�1��`O����]H�w��O�P��ˑ�J_?�� O���^������jI\&-����g�~ܪ��ՂH6!��WD
rۓ�}Aʳޯq��B0�6��C���
OU��r���Tڍ�eWi��87�4�nY��= i��Aw�qJ��>�4ȩ�q���Vs�"�'�m��~s�X(_w�>��TjEo�!�f;l��l]��rW��~��Y�|T���0���~$)B]�$�/�;������=�����=���mo-�c�d��0�` �g�
i� �L�{w��+_��6�͐�?�|�OK3�B"��z
�L�|��ve݋y�I�Cj�Fj�������oP�CeMY8��h�ڈq��tNw�F\aK6��q�����P\��{�k��{�����$ӻS�xT�BQT������B����b���E����5T��f�:9�n��@GIF0�RGz��"��[9�����X �Ey#�Ε��dc]WA�>�]P�Ի̉nUИ�fB��̛)6����sJ�C�I֧�8��<�Güdt���'�kI�Jy��
�O0���ۙ��Ҟ�Hw����={6�q������F��T�A>��0���X��p�'�r��k��۩�x0�Uѻ�3bd7�~!��H�R�^>'ӫ���%�pPh��X���`�U���������QV��xӈ) �$8o�ՀdZ�;�%��j���x@�O�A�(�`��4UP��h�z�7q��[į���Q� 7,�����c�:ݩA�wzK���o��/�po!�%�{�t�'��̗~-�ΰP��ߎC:P7I��F��d'�����=e}7ko�K�m����bD�zka�+&�dO*�ȣ��B��.�E
���M�	OX�K�ؤ�X��1��K�a�7�e
��f4/<�+7M?�=:✵;N�z"V�4+xe��&��T�B�@_x��E��H�^�lv�o6�Z�+��w�M:�>"k%r:���ՙ��y9 ��c��J�<OP��θs[2O��R#s�5=cv|��	�zMܹn���F/�ƈ�)��th "�F� ���LvP� ��h��<��Af;����K�I;G�����wv�s���)*]��N9��ܸUjoM𥹅h����p��!\�ڌ{n�۴F=ڒ%�P��0�*`qm\�m����XƳ{�:�5�EV�=������Y�s�!~�j)% [� ���6D\w��X�nN�E6� b>���y&I@���(�Z�*�gI��w`<i 2�YZ�X6�>#�b���2�T$��/�����pcE�?8 ��6�qT
�;�N�Ih������6r0��و<K��� G'�r���]f%�؆E4᜼�8�:�oX����O�Ĭ
�m{5,y�j��Dh
H�Q�j���VJ�я)wU���T���W�H?¬���K>)����Қ}��і	qi,��q����=ޘ�=Fw���LW�
��"+e�p���S2k��Thȱ������f�(���CBZ��DU���1Mb�Vd�yu�ל'�Xj�_�'��o[ej�p�@�e�?1�]6W�����3�=l���+%��Ӥׄ>c�I��+���r������_n���1<>��r�?!x�M"es�L�<Z�S���A
"��P��׹�J�Es@����V'aq��f^|�>�1`�/��¢}�V9k�9C׍q>�r#Ze�v�au0.#J<��*xI�:�.�B_��-�A;Y�Wx�T%� iB)1_L��+�%��\����ORr,b55�9i[�aȐ��v�{=]�n_mi�sV�kc�ypi��w↔��M�I��f��3��uƎsٲ�{++��P�K�+��	^]�(e�؝���@���Ȅ\�WKճ�n��(�q1�r�7Nb��j6�w���K�Q�08~\�����3�J0��,ش#���j�Ԅ\|�����лkt�;i{�
'��2���D�Ǭ^f_�W�9�E�'=B�C��M�!��
�R!��ݓ���(���3�v7�!��ח#@X��7��(ccmr+L�?"w��v&�P@�5"H�ݳ&2��G4O�y�"���h�2?=pZ��w��@�`\ذ�7|���#�1}t�4��eT����\��@P ����C\�G�d�tvI�`K��_#��RCE ������+�+�İFY*�I^-_^f=
g��qn��c��<~%�+��@ݭ���ޖ�j���0z聩��BpGe���m�>P�
y�[�!��j��hU�c���Lշ�$'�2�k�j/Lμ����D��R;��+Qޟ�|ɵ�BC�6��k�9\z��YM�����1�0��Qʇ�������P����C*����(�?Y��w��h�z�W�C@k�<t�e���^����>��];�_y�>���z�VXA
�8{�uWTq$��̀�&�Ćr�r���m�_t���#�;����T�u�H~���R������4H���T)�s�]�W�Dաr3�{br:b׋�k�n�ʐOD��	V��!�.`0������ف�݃N3��t6����li���1�{���.����S9 l�)I2%�ƺ���N,��#EE����9�D(��=u65� =8�#�-�/��v��R�gĤ���r�Y�BO���Y��-�,���X��	�Q2��: ]�oF'����9�U۾%h�Q6^;&�KN ��+5v(�y̲+ez�U���L)4����O�6yƑy��K�Ls �<z�KxU?H�2QD)h�f����v�Ύ��ɴ�%'�����u˓��f��gܿÑ[�)�^dʯ*m�����إ����V�a�ҥQĐ%V�Br�+0!�#�s�u����fb"0��6ok�SC�,��@��-z��A�ǦJ}p��A�-�ǀƇ?��·��܉n�]����k���s����衤~D~o��������p\�������R~vWr�(��A��N-�[���}�A �\"�����]a�_���	֏���C��.٣��T��࿣kY���߯��H/$�Heڍ���� ��/)�Hg5���$5GKiUV�X����u�ou�n�᭩�2<jX�;�\��3�7»7>M0	��[ʗ�Rz4���GG������_��ܨ0�AP���H�iUvy��0Y����G���֢+�B;���Yx�s�c^�X��� dd6'�[ZH�����l�R�D�A���m���0�Iz��F�E�*����Ъ�� oZ�Mf�ߏ�۷M�(�;U�k/2�t�P(WoT�l��5BV����:{9��$@,j���a�Fvb�0�C%skPbR�}��%��{Ǖ�L����.���5I���g��M�e@�ԍ�wr��1�#$�OCӱbDr9Ǉ���J���N�G8�)ܤV��=�u�9N�΋hM'�nlm
ܾ���8���䐜}aI�A@��aP�������d�n�CH�'	ⳣz��A��$�C��m���7�����%�{��Tf@�y�?�Hw3�l�mERap´�Q�A��[C��rP��&��H�ȵ�f��uӻ���8Rѱ����.��&̄��\�d3�t���N3�6�GP����,;��6����vz�S�i���XUd����j�%��G�i�Ѣ0�P�d�G�Gf�ԏ�\�����A� z��94�yҴ|����H��Y�48��
n��v����~��\o]6���[K}� &�j*���T�A�ek�m�(2���RBUЮ�(���Ϭ������	hC?���6i�c�n�((��¯p���"���[#�U��,�|ܟY0=�=63�Fؒt��;Kc��h)j!d�c�KC{���
6p�˃� EfPa-�:�&*�iZ�;/<�@�g㫋���?&8�!j7a%݌O��\yo\�=����5���=�>�Z�B�����̏�D��oK�k@�e�Z��+{�C�'������.��@8zW���j�����>&Ny�%�͇�rְqHu�@�41Ņ8@��AI���_ػmUm���x�>J���#Q޽�V���1��~m(r� �P�=|ip�`B�z��炴��=�Dm-�"�+�̹z��8ʙ�G..܈+�h��F�G�����M�ay��T<��m�s[퓽����`�]$�����/4��;R��݇1���*��-{׸C&��6�sK�M1q:� ��iQ^)ژ� fٌ t��!�.�r����@0��
��MUE���[짹��z�A	��,��&;��
B�d�WMx`ޅV���,:�>D���������&��_����L����r+*�mcҷ��/�D��*.�S�yF����
��dp%�zz����B�ҧ��h-�>��TG��_���;��������Ju�y�B$;ғ�"�Ӎo����3?��+_�+��Q�\D�e�چY+�Y�G��o�������Ӆs�Ƅ�Z��/$8o'����Ue�[�A�PWq�3"�Q�n�����sM�?�Ϙ�œ�5+gO9��W��C���q{-VP�o{��[
��鸉_��6 u$$Ӊz���.��b����cL�^P��	�7'+^�l+������;���7���A*�V6�$��~��V�����c�~�`߈i\Ȉ��;U|~F0��A��F��������p��A�Sp)aeW�Z�3�!+����&���	?�i��c�s�^:}-a�@�|A��S�}n�j_�(�=ID�	V�Jk]"�2Vv�6'K �W^ȦA��u&waF�������׃�R�.��ڛ�"��l����\��Y"�C/MYU�G�+w�=]|����f�-�SS��E��hg`8���b���!ܡ{E�L:o���g��r �h�9s�X���(JY"����i��i',qЦzeGi����J���A�e�.=Yҋ��u	NS�˄PX�1=�Fǉ
�9���4��6P�F�0�:�(��q�N�X!7�m|@Nc-*�q<����˖���I3��� �_�	5�h��FXD��7��ijkC�+��}�u���  ��R�!%�O�n�Ҫ���$m����Gɹ+�l�1���F1\����!e������?5�E}(ne,ɯ���ilkpa>�v5��=F�K��zu�.�:,[Fu�v'�6�ID��4ׄ�)T9Ϲ�����dC ;�Pޖ��ϸvV�o���/-�5>�n���Ё�t��H�^��0өqQ��$�a�w�N�$�K�'<g|Q3{{y��k��)MFg�P��	��ӡ廩��,�؉�=h��k,�#��!+Ŀ�V@Ƶ��z{*f�X�UgjQ�N���㎩d]�λ7_1�/D����IPf�!�3NjU���o���z�f��m4!+S�����C��J�FCY1ɀ��p����ɑ��P�	������^$�SN�X{��Y�B�<�ߺ!�0PW�y�\F��n/��IO^z�	�%���0��GSnj~%"������1�^}���ϛ�}����ޝU�8������3�$ �Q�K�k��M���ʅ^�����K��b�ɕٖ����ܿXM�УaU��~�@m������Jw)#m�N��L2 b
������UPMrR�V�l
x.M۽�=�	��QHr�]��b*_o4�׎��K�=�b���Q얒/����RO�dǒ3ʢ�ڨW���0�O�����f6��an` p(:�C�6�9�vh#��t4�3G�][���S�#�yo�`�w������1?�]�ή��b넠L��j��
l��E���"̧.�3S�EUCנ��-��E��rP��hs�G���
����-�@�a6��Q��l�F�ɭ�:�
?Z���A/9{/�Þ��!��gz�\<Hu%��[�r!�S�� 1��x6B.�{^��RG�����x�A�z ���LzIg���u
uM.���4ږE��W�x7ྸ.!@�$j�|�2'J`^b'��u�t��y$c��2�l�9
:O����� Ȯ�ש0 !�4����(���q�x�2t�4�X�_��������oS�;~ڥ�.Hճ~C�r��=�j双T�)<����	apIO���~�����(C��7ݛ�b�%��l}?=����OX�)ؗf���4HK�@�>�,m�5\ۃ�G�lK�@�b�r��M����v���l4�+Iz(������y�P�@$CQ<�gm�āC5++2��7�@�)=Dd\��ۃ0U{�A�?7UY�E^9l�aE#�yi�y��������g�Hp��vn�Y쀃��y�^*��Ψ����m�����p��@�A,�<D�qI?�L�ȝ�0|=�N�������.��i�=i&�/��M�O����2d�4���$�y[OK/ۂQ��C�����U����`�g3KZ�ш\���bꠢI.�S��Z��{.�sRh�3�#ؚ�m��>:��4[\Z�|}5�D�ws��9��g��-(�FD�;�Ƹ�	ʘ�=��Z�K<l�Fi�b�����>�W#����>�]�4��5�K
Wg��8Ad�R&�K����:u����`F�T�RY~�Tv��ǁ;!R�L��/WVݵ�6���R&.��
A������|y�v��'2҄���P�B	����.�]I�_���"2�+�k2���.�����n�1ޡ	+�l7��Cܑ΢�i�������e��w�I�ˠ�Rs�u�֦��Z�򱹣m֞�h�eb� ӌrWYa����$�'Dy� �����a�x�#�]�����FV���p&3bԳ0�	2y,=����3�	s�Gr�(���y��$������<����X^�bak]�),8}LX<n}��_��|���T�O<���9޸���@z)�C��6H~r�5��`"ԩ�|N��K�9��<��o��WM�֫����}5:W�;���by�Ӟ�k��l4O������/d~��{�����ؖTRWN\����������#���)�0N�x62�F��K=E���+aRPD�"нb��^�yB��ɛ!����$�<���S\žv���{��n�������� �_�	�O��isQ���q��Sß�mS��;zթ�����"�1.{ag�S�1/^ۢ(�ߺ�y`
�m�[�dZ@-ғ��@�c�̈)bi���W�-�U��ew�B�?_��ŴۆG�����y�n�����h�/-oq����#�
�2~UU+���!*�Vd���͵Ly9~�ՇGs'4�`�!| B'����I�G嫹��*�,i�]��8�r�l.�:#���=�e��ꏕ�BѦΝ�z�l +���>�r��KOTWuw���	xJ-#��Y&Z>�C�2�2����-,��T�8q�<�)5~S&ˢ�\�.�PfZQ]υ�,��\l��Ϟ.C�D\���T#�G��@n����d�	Q�� 1���q6��򒪽��i54x�ەg��o�j��9	1/'M0t^:b�գ\D��.�L>�`��T�,���J��0׉kvg�� !�je�B�>�����XK�Vn��7��"%��xQ -ݦ�,�A�>�p���Pn�O	�:�k��b�cg�}s�$��J�?�M���d�� ʯ3��-�S��FXl�� �}��ĵ�Y�d���X��c� ���~; 3��\�PsK/̮M����,��`�p*)��W5@D�q��cN��v�4�I���N�/ۆN�}\�l2K���&{#�@���W}"C�t���t�1"2���>L��o��8�Iی�i4KǗ�3̻P�2�d���8N�$B?Mú/��j ���J��U���H��I�Cx-� ��VI�w)ѧwuc�;4�8Z�m��v�j��(�d����~g/�(��` ���ڿE��j̛73�N��J �@�,�QZ�-���UIt2Qm��\���b��%���C:+�"ұR!@���n��k׊֯Q�IK� ����bKU$������U���bٹ�����WT�L6��}u�2Fh���Ej�r�%���N�>���I��aWaJ6=�y�� �� �Q�]����Y���u{B$\R�/q���Dv���1VYL�j%���,��qR�u�Z��HIOW�&ܻ�i~)���FnV<�k�]V$��.1�l�'iH^3z����4]�r�����{�`1 1����:k�p7T���tt#?G5�$|^wV����	BpKI��$dx��6�;$'�_�G2<� �t�1�2!S�����~ꙺTR񣻖����9���NX�Q����R.� �^�����^bd���j��BsJ�ܵ	Β���mT'-�#�Nb��o����8��ٟ=pV�:j9w��221�W@�lB��*}�ᡄLڿ;��;m���$/#�yKB��������?���Usr� Rʙ���f�󾵇R�(:�'�T�m��ƌ_ƝS5�p��& �;��1���xu������q�?����q�nYl�ň��6�3F�
I�q������2�K�fQ����4聳FHx�]��������D�L!>uU�}���O�y'^� �G������o�h�� �$�V}�L�aX�:�k)�;.K����J�q�����2���W.K���޶�!�� �%��p&���m
�����{�mZt(�{�Rh[+�*�qeҚk�zW��1�#�iIC�>NM>��a�eMū ۍ���z����C��i0yY����o�w$� �	'͢&x�$�饵`<�<;���[��j�D���/�JY,sUx~�t��Y~�X��k�i5��)���NJ?�R�d�}.d�I;�J�n�	V)���]��J{�G��vV�)� �+��1+Gx쬾���8�P_�,҈4?i9*�N�&~/a�~�?����*���L"�W�R?d�hrz �����S���XȂ���	���M|/Ȑϖ��ɑ�P3	�L�Ma�#J�Q^n����YӨT�AVcJ�>r�)$���{��X%�J��#�ӡ�v%�ղ�}JtVB	W.8޶�*�D��-���P�}���94�SL��!�叜kԍ�i�sJ�����=��Lu���pnA�-��o�-w[��=e�����a��e���lc����(Ut��A�_��4�F�sä�j��!l��	�5�`�>�S�5s{^% z���������Q>ڌ=��"	|N�,4+�@;����J��l�KJo�.��'��jܛ�Y�}�q�����:t79c�ļ!��A6L��K�r�H�k�$�ѡ�2��=Õ~Z�4�[
�0�
L����N������,7�;q!`Y��g�):�"�J GD�r2n�2CT����Կ����xe	���y�kİ�	 e���328p��t��g|�Ǯ�[_�N�3ƿN�GF#S\�������qC�]+�	��=U��=84��8��/a���0Dg�oH;�����W.��/�K��$~�V��۟b튣�㌴s6M�av��0���|n�B~&�ƪ����d��Å~�Ս=Hs���G�m�x�~����g�m;G��r����H6K��?�2O�;���)J�5��` 1���.$�c�2)��L���*���i�G��o�6�x6��M�6آK�5M'%^b�	��4�G���a�&�;H���$� �����Y�-h�?�7��h�����8[�V�g�'*�s{��p�\]-)�-�?��\��X��㨒}Bzi�Z��$��ۙ E�r��iܚ�����=���]|p�=J�v�e�`c�y����=� P�7",Bߤ��}��W#�������,����/2��;�,!�F�c4`?ڬB����Q×���ln�6^�����JU}l�Ȥ�hE���t�*��ǯ��g�?��La�!$v@}��DA��{<y��P{@�V%*�����1w;��2I/@֍{�L�g7q��v�A�e���k�F��}�Y��y7+0`^��A>��.��Y�p������,i5W)�숈	�H~o�~�̏������+4qu��gx�/O|�g��x�U���(�v�A�g܉�z�}Ӕ՞�&�<���_�?8�n��%�)ܙ��ƨ����7h�'ts����V���V�t	�O�'?C����]���1@GtKg��\��f-��)7Go�^xy9�؂���˽��퍋���\�՞@ʇ��7�.=�GO.�e|G�NA���X� �R�+�|6��J(v���~qO��)��n�x����FU�d5o@�i�ʞ�E6����dK��P��a��i������ ��z� �*"��7� Q�`	�sZ��.���� _�#M�x$�=Dd�J��!��ZtJ�UU=g��c�E�j�yҊD�fV��[-k��"�������F����dL�";��R��ߍ3��ʍKRRѪ <�w�ԛpp�x?0lL��:�e��V�
�{���!I�N��~$;-��C�x����i�3vjX��h���Hˡ����o��Wv�|a��t2�S6C��A|x�e�B�7�R6uj��1��̬��̾(�u&�>y�Y��XH�a��+����1Z�?�g�1�k6]X��$V٬�N�E5U4�^�ݥ=�B
bPt�@����d�t�+T4�2��'P��ó��䨤��5s�T���d���+[�^Bw��wة�|^�<�U��9ɟj2P�Đ�t�O`��N`�N���cX���J�M�%�+�T:��?D:O�8�h	���j�2�o#}��U��0����e�kB!�D�'�r�l��A1q�RГL%v�\H��l�2!vO��);f����ș�tH�OҼ_��$���c�8 �\�Sͫ��Q��RJ6�;[�;u|54�	�]å�f �~����r1�>F��d�|���EH�G��.��/���|=��w���6�Mn��P��;4�^�5~��	NcjD7f�Q��w;/�bdC��d0�JG4���V~�A��,v���ڷ������<O�T�#5:^�֟��m.�
]�p���W�P����a��M	]>у��"�b��p���11̮"δ SU&��*B�YHxEWw�.C����J�J���1l1�|3��?!��3���߷�:�0��u5�� �3��KvL�]�?*&�	��\Ȉ�6�G�;5���ſ�:o#?�-9b�i8%��/B�ӡO[OF�ME��=�������a�X�a��{�ǯyA�9�sN� st9o�Ll���H-\����R;�r��s,5a��Ơ$��￧�Y�bK�ƾ�ҲlI�y)�*��U�,��_P��أ=Z�/�E\Q�l�Ǿ��@1�t4%Z�S�V�>!v�$��04oF����ƴ)N�e�g�_\�t�U�'�<����t��G�>��7��I�k�Wy�J��藚�/����FP�_��z��s�oa[vԶ�Sgu�����U/<�kj��>$u$@��EL~RH�x�(��n� /D�tͿ.�eX��[�Y�H%�>wQ�B~�h�%7<t=�M�;�_��I>I�A��b�������p�|iR�jE�%n4��[�߷�I���P����D/>���G�6-��v���O�EA#^q�����#�r�a���!����&�}��a'M��r����D����Ss�7�U.�]jɯ����ȯ*�w|t�'eu�(��}e�ơP���m9���Kpis��7m��'Bw���iO���|b��3p+���݃Zm��{������E\7�?���Y,d�~����`���˟G�7�*/hۗ�v��`S�����T�;�����{�FŧK�y����Rk�[��ꉹ 	�gv��Gc�ʝ�d������R�et����A�!�"�f��?�;��B�>k�S��z�.��{���C�#��v�I���l���L���2���)ИwfT��q�PXT�����zݣ�S�W���k� �ЋI����"�q�v���\!�R�r]2-�3H�k\�d@[�<����!�g�p��L7���x�A��/�w�d��9V����z�5�І"t�,����f����t���1'���mFE/V�㦘n�>[�/���50���2sЀ��X��6[���񮌘�}������>��v$�M\���CKt�ْr�,�����ʷ��E.����!cm�|H-V/8�ޝ�0�3�k�I�9s�%Z9�J�6L�~D`�6:����7%�d@��z��������%�'V��*���3'��P���]rq��H�i��P�/ƧD?:�3�.�J��N��{��i:VIs�<�$Z?�%3��i�~P���O6�U0Z���@�����m�.38�$�M 4�7\���rR��-<%R��K�"@���[�AІ��L%og�?g��MFo҅oX�"-���Z$��KP)�Q��`���D+6�^��M< r��	T7��<����g����R��^��\�5H������`A����� �޻�?��Q�~aB�]`���*(\4�Y�ܡ-x'�@jgr�B/pp�o��qE�Y�����U�W��=��^m�ߦp���r�0�IL�2��12�y
5��YuI�5�oN¨�<�m1��Nn�uN�J3����(�Ě��&����UZ�]Sn�\����A�����Єr����"�?(RZ�H�����y������T�`�bPŐ�a�j�����=g�O��1C����`E���8�ڲ�y.���sGH��8�����pWe�oFT�m�cK�!-uͺ��p�p��=V6`�5�����������y�zl%�:Q��XQ����g��p�?��_�p�$ٜO`�<�&Bz��`�n������r^��cb��NJ�	德\��*l��j5����x�: ������cܠh
�~!�׬�#?��g��U&uy�l2&mP�S�;wuʞ˄?-���/�����W���(Fv��ZG%��.@J�_�̇�QulX��7�~_��%�ˆkq+��bF�H���-n7�jǮMk+Q)�`���}�2{`F:�躎iNoU�g���.�R=�H�g)�5{���KzYo-��m�->ta��Ϫ�U��H��I�oX1tD��e��u�( ��&w�-�n�i >n��R�-�\�k��Ɓ?ef������gJ�Q��	�$l���L(��jz��_�kg�{1���T����#�ҊD�#�Y�6ȵ?������Bw���'[&�?TҊ|��'0H�q��O�-;���5{-ۧ��1��|�n�Du^p�h��Yk�$�������e�H	��^A}E��ZP�v�?�M�N��T�"�����$��5]��`�Ȑo
MqN�x��Q{-n?��W�L��:�:�J�����H?A��|E�q��<�<��+h�������cD��ok)դS�Pd�>>���7��WGw����*cL���!-.�5A�y�e6���FH��ʰڔ�%_$!K���ÌcW��&E��:�7�C��|�FjӈK�EX�ᠺ�d���%	�*�R�I��_A=�#���<���,�6�,�َ^R󪨪�"���gM��+X�=,�_�"� �o�����Kq��d���d^��]o�&�X��A��c4���A�n6�����~_$?�5@��6�PF ��j�դ\�䤁��@�|��DN�B8�FP�A���`��~`+|f%��di�h�Xٜ'�$M��Z�,\��ƴ��a�/�^��e���럍0��)9���۸��VҋWi���j��e�����`�a�O9P �xr�+�d�E�K��Q�Y�N��j2k�*�[#��of[�Y���X�
�_�Q�FՈ�T])��SK�������6���7x%���w�h3�������������i�II8vLi}�x{�cvq�"v=�܈��%t��o���qi���G�7�]7l�q�6�&��ˊZO�Sq�.����P���z'Ҹ���򝲷�*N�oA+���%����e�iX$4#~1d�-�LhYj3ـ.c]���HvS��B�Cc�*7�"\����e����S���ZT]&��8w�P�.%�{��$k�t����Hu�#Jh�1\�a��?O�aJ�w����k�M�(:�JX���.��|A���$�XCS�#�_$m�4�H^�W��O�]j��4����
���E��q�1��7��Zp��!�K{c��x����]�����R���[�CP��в۷�c���P�4#��U_>��)�>��S[�˓Ǳ%i7qevH#�W���������&�_�S���K:3�GB�K���Ay��[rT�*�/�<pG,5��\gvc��*8+z<�XY��Y�6�Ic�Jj��5V��������0�zP�+Zy�J]1���^�q�����d3�}k}��\�㢭�,��P�2��5Y�V���zF����%����&@�ě�~/���l�Q��n7�sΝʖ�c ����j��@��h��"�N�G����#ҽ�.�V`��:ܷ:o����\�J4ﱨ�
B{�·��~��&p�3<M��``�(P��PMCu�Ш��B��o9ý���D���~�F�� ��Y(5�~2�g��;Ϲ�P�9�ӰWXY���=�%��76 *����k��o}��^��#���L�E.��䇽x��è�3�˳��w��2���S�=�����A��,lx�%�����
�2u��E7���[��~�붶I�0&6�n$U�ޗe�/�;ݱ'\��%x�,�` k�!:�� ;��H�A����Է�����YCh�N;�~LP�v�0�����J�}ڛ_�A�5?``A}��'Xj��VR��=��S7��� ��9�yw@�sIUID/�6��>}>��u�ȭ)��o�x��eQ�d�����W�6������=�}yMC�$�|KӸvҍ�y��f�QIb;Xfuz�:!�Z+�%��DI�Z=�M§?�&�.���Mx�܌ԉr`��U�{��_'�*�и�Dv��V߁,��"nq��j�zo��n�(�N��_���|�z��;s����Uxy'�5֜SWzSu�����H#��8>g(S	]G\A6K\�#��=	�
��ᦅ���e��/�a���=����S<�=}p�JI)��`��XEzc藞W˖U�>�Y(�EԖq�W�4+`�΀���qVO�Au��~,q����%�J��W�|�*S��O�ާ����v���G�v;B�=���e;4��H�����*�����Ӂ��㇙d���Pz��x�� �ߧ]����̊New�Y=,��
x���J���ٿջx��tO���ef֣��x��)�p���­\��)�Y��=�8ɴ�IPA�2�[Ő�?.l�m��� H�}�������8��q�%(��x֨xOws0z�򶑆�X q��Y�PYC��P��=����0�+��Yi�?B\����������n����K����wT����>�%J3Rt�D��\P��F���ԋf�G<�nW�4��{��5��h���9
�1����X"�&M^^�:6QM;����c0�9�c�K��q��A��(k�<�����g$�gc��#0aJ<|x)I%�~K�M
/� �]�
[�T�!GL��mL��6���<4�#�ͦ5�M$���L��#�{����g܏*r%Tƚ��s.�H��2���e�|�Z��pci�2 RZ�k�,��9������ߴ�ů�%u ���XNk�`�Ƌ�qQU���|��ΐ;�)X�SO�kK皆Ro�Q��Xk�UE3h��f�����2�������M�2:DL�9��\����������/�N��9i��>�G������"26%�q��ؿh��y�f�Rz ��(�p#��,�z��I�<>��{S����/��B�/�N��%�F�����	�,��5��
��.	d;]�9-���=�t*��}����W�;�+,&��bU����jV�NcӦ� ����]��|Z`[u��C��<vWO��<t]�g!�_Ԣ2	��������ru�j�7�e'!P�� ��?@R.wg�j�r�4� Ve�Y�e�Ͼ��rHo�3)���ӁDq��DCdO���k|Sx1�q�A�7 9��0����#sɻ	5�����g$Ż��X�d��օ"�*����r���wՕj�oů����x�'!�V���(=�evQ�5�/�:��F�W_\���n�\,^GB�ޭd�F�����xڮ�6p]�>��^0GW�j�x{KB�嵏�n�*���j��9�g�&�������J�_�	�M�Aj�E�5�>���������	�SؓԱw�[ci��ə�w]��/��׶�C���`$��ٗu٬����"Zѿ�����G2���!9�����ㅁ� ս PZ%�!�_;'��2�Dk�OO�kTBGE�����$U�oΩs�3z��h�C^�ӹ����G�E�S$��?��o����x^�{C�|T}�G�B�tH�7��a,��Qf����―�442�e��d���M���@f`���8��(�\��j�Up491@��|�A�R�W^�g�t��^d���� ��8�l&��>���7^��mK]>M��c�r�p�C��=�R� �d-뎊���l.a����#��	��nS8Ћ,?�Á�Y떯�HuG���)��|�L�heI�l���4��
3�֬��HtAoXZ�� U��ls;ƽ>
zi�л�=�� �V�>�`�j��3��d��4i�p��ΧMrߚ0t2����|s�F��v@ל�;l������������*�;��]԰p��G��S��C����((�h�M� e���<�^��&�+� a	�	�$����[��'��^�?�}i������p_�;퉏`���dWB-�@�KmLF;�$�<�k��ΐڧ�Q�KIH�n���_Ɠ�I$(yY��ҕ�����nea�F��AvY����y_ q�&������C��$�M���1����u��9����<�f��	k=�.w(�Đ�n'���/��bh��߉_���P���|i�;�3�D�FE=��TO�_�Ǫ��w�kރl������H.�9�g�Ӏ�|�>������
*};�=�oz_�'+���!k�J8�0�
!�x�G�w��X�.��+�$�U��c����6�}��&g�:lMv���#��NDq����1p.wB�c,�ޑ���fȥ����uH4bh�O��o�~��Uӣ�S��97y@�os]���x���1��Z�Q�E ��V@�#��4�h�wr纮yO��B��'��v�V�5�o���3&�I�l5���K��[莁^W���d��0/�;�\]Dv\�3�w��*htRN�)�4*T�2���?�dJ�����7�Z()�R�B��n<d6�tdB+�$�z�]��N�W��j�FP"���ywv��fv.��n��Y��SV>!�BMK��l�@��72e2mf��\�7��� T��'�B��riu��ؐk����Ur�
8���~3�O콂��֝�^Hy5ӌIj]�>a>bV�[oW��;�K�#gP8���*�a��X�N+c�wyXP\�.WV^TL�W"��$��ZZ䀱����d@��(@`�c��@�%��,�a
�����'��p��RA��U�v���9�"��?�(Z�/����T59s0��?&��-���8�ܛ��l�Os��O�2�bwjoO�+i��7xXc�2��H�9(-�n��l���u�M~��ր�i�����%o�c�b�zs�/)�	�@p����Ϸ�w�p�gt�����.��V���>�D�(�m߬��3�A�A�F�}�ѹ����*�7Y��D�5̴��gD! �Q�(�v��S�Aė�Y�K��n%�p2�?���5��l���j|�b� D�GB&�=@��"P�掰B�,���!X�Zj)�9�Q�K|�a�ذL�ya���r7��P�hTp� Q��r�(�p�OȸI#�U�)I�����-��I �a
#���!��G�Q��T�e�D��G>��t�uи�c�J�	��a����A��P4����}ll�0u$8���+��������Z�Mآd��m��y!x�1������u݁��E�D�E��m���_tT.;��vR�i�%١�72AD����Β>iT���_wXs�����EÈ��@�)��-�~�鞴,r�"��6֢�����8Ɣ�]���*�Z^;�ւ��`,�'
<+"y�dEW���>x�`�k�������{qۦ��3a@n����c�=����&�����0 �F��!,�}����5��h�y�-J)2��{\�����M�>IqQ[���4ϟ�d�B���Y�ap:ڒ��X�$�-y��2+�?,p��|9G";�A�)��wn�fp���[���?����kGC~��0��F��+��	Nk8�u�t����!�6A������,AR����sxfm�c��(���DOZ_3�M:]5\Jf�p& n�@�"�b�S���h�v-A��UJ��?�ܜ%BmH8�д��L:qu�����?{
�;����2� :��P�V4���u߬�a���Q��W]v��j���#����RC�Xv�d�~���ԋ$m<�C�dl��B�.i��gRI���5��Jq.�}���"Y�z�TpϨO�2�s�^�TA*䓍J��X�K5��N�`W�
"eI Ƴ���A���IG0�ᛃgA�</sj��l�Ms��v/i<u�li]�����O��oQ]���M��������ҎA������}�]~꺆�6�|&��>8�z<a.t�T�����]�BW����Mm)'Oł6����hVЋD],�M�;�ƞ�v���Q{׆���t��? �Y��2y�E����,�l�u>
��Rd��8/s��-x��D���a��%<��Е��c	����ԇV���ŘV���<�B;��/7��
���V<��[�Z���Ht���X2�S�_��l�7��^rO���ԑ�$L���S��.��A����W/��u��G0ˍ�K����	�7�m^���	ٶ�[wC@�����Nb�$5C�(�bqh��n)>�O��S����X$8��˒7����d�TW�Mn��e��'y44����Qyԍv� �Ԭ�'��]��(�j0e�ꌬ+�h�䤸$�09�N��y�./������JY�1Zn'��ut�'���O�pr�BD&����B�.�Tx�<۶ђn$+�>x���V���H�`�Yn'|��-)IDG�K�(c@
��)K�~�F��h�A�n�\���J��h�f8`�ogϲ��i!�!nY�0Pd��ZT�܉����Ŗ:��Ɨ����L_MˊX�}7�<�"�s۹@�lzs颷���f�����`�p��lw� ��E4n����>0�nf�n�l|.�eZK�n��&L������Z�i�N��Y��Hb�xa�*E����O䐰6f�U���{BRe��.ԡv87�%�\��C2���}2�泭��>XQŘU��O4_W�(�}�w'kA'|b�PP�~!&��*Bw�%�&};�]6��J�	�S7��Ո�Â�*�C'^]9�������s̗M��^��"��_��z
�5�֔t.���n�eQ���C�o#������H7j�Q�������n+�IX��~=`�M�����q���2�����A�2���1�P�<�m !�}0�3"���(ȵCwۖd�'�:���ή\�wnw�V?&�X���1S&!�	���f���S����>���v=��1��3�o�AV��o~ �$��ꢂ�[����c����:ೲ��V��� a�YG�� ��i�n�9g3���c��j+T�:QB�oQ_�=H�̄y*��r��M��Na�p��f���|������6Y�chr����'��2b���vʑ�mi���+�	������,�!�ǋdes�p�g�L�*h��X�Y�I􌶲N�Y��A%?��<v��������;�ˋ�$�j;Ռ)��F,�yl����������l,f��_X���Ǘ�c�!EP�NSq�u/A��v�:�F�x�9���p`�1�g��n���fFn�x�O��k뗅�RPOo" ����/�p�:�y5ǹ�&@E_<��<���@��}�9cp�+�m67�?9�d�/)7l<s�B6�Lʢ����>�Y��� �P%6�z�����2]ヿ�!◝	5����a�5�)�/�ǈXh�	]�
7~ �.ؽX��
[ }�����~���_=ӠT�kh9*PcV��K���=Llh��H��cX, ͘D��^5����p�<�O�w�ř]B!*����3V�a&2я�'��mwҖV��8�<��:��-!k_�M��(�,�qh# ��zT�q�����#K��7�x�8����2]�L�b\���8�PWg�üw:Vͽ��z���tc�E �bp�+�	�JkoO����z��\�=1vMirU7eX���;��9Y	Q���r���|=��a�2�?h�G�P�|Q�����l ~X�X�Xa���d�>�����=��{8�m��A�h��H_%.sȨ���1 u�2*�����=��|t�����3�憹t��p�1��E�b
�t�@�����H�c�lǢ:�(8���BQ�sڕ5O#����_��6x=�Z�A���D_� ޜB��l6�WǓ	5@̇�]L�H��	�H����Xn��
�hj_�ik����B�V��'l��>�|4>�`ek������ꮠm���U��I�dLG_�ilE��O3RPn���(A"�b�|�-H�> �[�>Ӣ�����ߦ<��~ �?���ʨ5�=7���T�Rhw�ap����VK�^�`��{9�]���܎^�PȻ�ť6��&��S5��</4��T�����JU�Iv��ǯ�h�=��*�n(A]%��L�+��jΔʪP��s�tˆ�:d�\ Q���=�H]��rw�>�]AG�������
^T��;���st�8���v~�GoBh�:�¢��cY9�<��Y1��{��;�1��ʐ�#�Ylu �-k	�(_��gI�[8������1i�m��(�xS����Vo�Ԥ�ʨ��9$S�H=6k���;��� [/��´��Ym�Иg��Hh�\��ץ��; ��9�5�L��-��Ic��z����+ܦ����s<���Ш�o��0a&�����X���3���+f��H~�W�'�s�,I-��)� tBy�b.[8ӦUwLߘ��U��G�����*.�/���=��O�<����U���Cp� �:�E�rp#�W�r�%�=W���9zx1bP���5�i.�Y����x�1����J8�%00YNؑ؅]|���������Há.�G�pv�,�/�KU;t�u*�Te�o�Si����+�#�I"���-De{�nBT3L�]�x\�6�as�K������h��2c�Ĉ�M܁"���[�����l �}S`���~��(`�Y(���ّǆ�1���^��{��y
� Ҏ�u��>?C��+f>=p�-I��9Ij���͕s]�y�3��)�U��=��F]��˒��V��ܜ����R�Q��e �Ͽ��y�ι�Q���"����:���u���+���yK�>�ڠ)�ވҵ�}�I�-�W�9) ^ϧ�Fր�=F}���M_3cd&��6�p���Y�o_��#Ͱ���aϳnĺC��h:#j���[��^�����4k����0�����C6���4���)o�����$�3s�� Öd�<��pN����2o��"�<�v�%�$����]���X�ᮤ���bG��uc�M�.��U����޼�u�w?@7f�A�oZ`�+jg�xsMW�S�:6%����?�'�(����ET�.?�	������n�e��I�����/�l�ж/Hm!�~���a�����n�u���*A��٠d��sQ��'�+?I�ܧd2vZ^��d�%��H�f-���#�S��g���s}#CL�YRg����f��ӊ��G���FIPY9&�!��b��Aܮ�ʦ�!�s���w��.�#gL9%W�������3�	u9��ĤC>����t�_��-e�yQ�j/��&/�-�M�L�{���}�V����\�K%=��9���~֨��A�\����Hq�q8{��@���xWV�a
B.��!(�������yD�'��R#_��<��O�%tN{ww�2^2~���
��^ěUi7.g����E��1w~�)
���:�݆ҍ��q8��M���~&N���#P|U�ϰ�����,q�����j|z�hu���xH`u��A[�B��Ȋ5Mj��ȇ�}�=:��	kE��Mc�|}���������Y��Ԇ:7��#���%p�O���!P�O��Z龷 ��{ }����Ȗ�4��`?H;7�jx{�[��-�&D�RX��Ⱦ�4�27���/����f��$m\���B/
T�x1?�P����
�D^{�+.uq�2H��+�tʬ�Rе�	���\P<[bu�_
�%��Zsf����h�mԚ�Y�Flr"S�����s���+kw�\&��-tFܒ��C�G�|�q������Z�T��&������z�V�>�QWR��u��8�W,ؖuP=,j�ZOsD#G���ӏr>b��|M��h=����wf�^S2'�>�F�����z���"��׻��{K��ѽ�l񹡻����|�M#�c*[˂ZdFJ���}���Ķ�LϦ�\G�1���)y�:)�Qy�����88|z?��y����z��Ү���c޽[��:���d�֪�=���<=��L�m�{2D���h�+�����B��v���u��4j�[Ժ�ٰ�D���e����g�/y����䭚��t��gO �L��n=�;�������t~�-R�=�i�\j1g��%���5�Fu�o@t0�]��ĳ�p�����<|=��X8�yʆ�̢+�xD��$�-s�	�a7����3'D��?�V�i�z{V��S��[����S�An�W�<3V�%}��G��������I_�s&��f�w�ە@u}�j��#�
�.��	^}�ջG����Om�j�C��7؎�ć�fZ5#q>��dH��!�6��y����k"���F��3I������(��=���VN-�7\�#Q�O��}�{T, �9��%���wu��?�:��.�@��}f�Oz��ו�/F�Ŕ�	[��jϣ

x!���I�)\Z�h|/TZ��I�������P&��G<,�Û��?퓞�����l?첥��7�����I#�=�Og�S�^�*4��_V��B���7'�<��d�����f�Y9����-�J�)��Q�u�~�n��s.����)�u ���Y4^O#5�D�4
��c݋g;.������tu��:�TܸG�Or��"� #���� 9΂ܣ&z-W�����dV�y,E�O_�?[#8O���o�Q����!��&�,zx�����~���D�[�8�
O�<���J��e1r�ф:	�����d�)aS�hia��@���l;%�����9�\_� T,ņ-��KO����m�C)�B���}%�|���5��Џ�c0!d˶I���%�S畧��˫3����_ �E��r���NWp�T�՘)}'FY���$�<
t-(6�QtE�!Bc��a S�A�U�9��̌�S��K���<��ˑ�#'� D�b����H=G~��ʒG�5e��u�K����^����Ȍ1u�S�L�s�Nп<M�Q:T�Ŋ�^ޔ�I+٤����@�̙���(W$�BC��E7}�Ճ�f�1��?���%�x��������X( �"4��e�@}T9�MV��`�����4��H1k�pv�.�X��3��V�/+o�:��4�v4whz/���z���'�w�S*�ٶ����x�ب����#.� (���^ ���7j�u)���#pM�����`�H���^W�3>Y����s�]���W�1�����<~��4�2^�l
�������A*:����M��o�)�d�#\��_��v����6��Z��z�:.0Rˇ4� ��G>�C�Y��0�sv wk(�\ؕ��??ult�8���{�L���L����bl���
F�WHK#�sWH�JS�����iO�Y>�^D�DE��Xy�&d+��,�g���Z��n����$.�e��KZ&T�b����*:Ɠ���ՌY�b��rө���xX�:��Vz�q�����%d���	�P���?�ƭś#n���;aA%��ֽ�< �d/�S%d�e����q���ƣ�A��
E��� ��aQ^%Eb���@c��TBR�bhfp\,bo�V�t��Ɉ��lCi����b~�J�N���^�rd�z}�{��)���b�k�IG��2O;.;Cj�7e h(�O�Z�j�����HM�n^�r�t���O����Ai<9����H�>-�FsHa��٧g������p�5�ρ�漵zP �7�aϪ�N��S̋E�oo�1�I����FNK�W��z�z�*��D~Qs���Ԃ�����+B
�j��F^ɯ�)�~���
��d���ک��uom/��*�i�=���\Y}��C�9�.���܊�^�"�|���c+/"�!�~C�|O6��V� Lj��'f`h(+h�Q
�ߔ(<Z�)������T��x3L���l��B�F����&(��ѵV�-��}0r���c�u����p1_����ߠ�eY��$��Xð�o�~:��NM�ӗϪ��cx�W6(w����XB>�ĥ,�U���u%i�G��)�w;�mTA�۽�q���ۨq7����ҡ�����r�G�F�u{����?���r�R�������a��^�D9]��u��6ʥ"���.Ao��Ny���t����d�&��o ���)�{�?����~V���[�읧[�K�ڪ�%��}�*8mbq�A��Y����`������qϣ��8'���?��;]l��U9��؈�W�z���u�#��?�_DfN�J	�sk�a���V��i�&����%!�b#&�oفO�����ia��]�d�TT�:w��H%g�tU�2��=|ѵ�0�w&ݱ'����>tOx����r�y�e'>r�oH�_�PW	�EY����'����Ŧw)���B?@l4W`��ȯ�>��nƖ�w�͂�$�>06���r G��<��e����s:N���j]d�$�9e�#��H�D� ĶR�d\�,�LK��J�v�'� �~�VE��
��Ua��6�\w(E�9p@���Q���K�!u�T�E����Y� ����AQ`��>O�j秸�MH �Uv�X�]6��nC�����������~�b*��D�ak�oף�l{�6�ݦ.�!|�ٶ�PM[3>_�浞�2����� ?
�o�+������n�<e��br��[�i�@�fX���ʮ)?FcV���1��K���0Եǹ�
�q�;S��@�3ut����HS�W}�q\�<��d54@@M&J��r��h^�ԃ1�W��\9B��j�	%l"�I�_�"W�7�7Ҕ��Ί���P(&��)��pwQ���%a�DF{�}SM�v�k1��t���/�`е�cw>�>?a�� �x�n��+m����n���J״�\�/w�d�a�$o�X��
��cP�o� 7O��3e�l<�è� ��Xܒ�B��~��b�K�S��5�'m�A�{}�(��<����i���r�M��1�K}�E�S�z��[���~/:A�K3D��)�����:]2�X+۾���Ξ��-�\U�@K_S:fl�/#��F�w-�ۑ����R��!��`t��`�6��<��XWS�Rʳ
'�&Bj��I�(8l���ok���%��<@υ}���V� Y: �������ܥ(�������6�1Ȁ+��~��i�k<7u�t�,�	+Q�������J=U�
�=JYv~���k��?�n`�j]�%��g������3f~c��#8
 �����>�q�4re"���8u�Z�'9U�)�#��+ţd��`��$��XӍ3u�D���������4+ݲlhL_DH��Z<�44�\/���R�ÂM�4wU�k��&!��Ɖ�W�F��h�j<=V�%��ǫ�HV��	Q�Zj� ����qI��}nJ��Rj-Do+� O�b)�������>�]�z[���Kv�=�V�Bw*Y����dUj�4�Q5'�j���A;��r��F�N͟�U��M�G�v�P�c�g0�8�pXZP\�"�\\$���츼k���Ca��x���jR.z��;�����-$�����Q�{z�e��e����|�&�H[E�mk�XT��GW=߁���c�����IM���뒋�6��;Du��[*W��@Z�����v�d BB���`$�I*�����;��%�.���g`C�LН�G�����������ا�L��Q��"����z�0G|��ٌ7da4������e&��H��-��0ܴy����[iŖ;u��A�l�_4�'�s���Z�uĦ����ag���/l�ҥ�.ބl����@#�����o�aj��+��H'��.���W\���6�����_D�;zC#~,^u��&CƲ:�36Q�A����j��	����(&qg;)�I)/�
\��V]�~=X���Uͬ(h�Hy,Y�}=�x�nԭ@����z����n�Qbt��LEG�sy</D�9rz3+�Ps9���~"_���c��C
?r�GJ(G�Mj~��*�VǮU�.�2)2��A�
����:=����=ֵ���"X����l<��*ex{l�Aօ�J��c�4å��%
��Sj�6���9]�JfW��	m�������|g�dy���D�6���T
�
�jk���C�;#ܿ�ї�ݜT�깵�4��t�J��^�r��"��}<��	�PM��_��P����y`u�f�ߔ���l]ň�h���" �:�M������J�)׺h�L[~z�x����P����eKǢ���E?͇/8����:��C�=e8f�� 3J$�S�gɝR~����ԕaF$~�J��R��rv�iĽYJ�
�a�MV0a�RO��r�R�
7���l�.�C�(b D��Ĩ�&�`�'�ЊyO�"Ig/��U��'��ه�[��R�2ȁ���qq�>�����-�c:��'}��wq��+����<t�0C̩�����T����3�����+^��uث~�Ğ�c��7�3�-�,9E���8^�癗�N��wZ�}��i�B�ǿа>�NX�byO1�+�L�ɝ�q��.I)DE�(�������t�yuag�bF����"C&.��C_��>(m���{�	3Եg*!|J~��.WW���F$W�u��[�8���N�X/Sq`�[����&J��۞�]��۲��0
YTbl�w�	<��V�R@��۠�#7�evԚfBd�2�b�ڭ�D�������j/�S�@5
��ئ��Sk��ޣ��\��/}nf�
F�!!B��?	X��0�`���������OjT{� ����g7���ΣL"?	P��c����R#*D���zdD퉞�T��:OE��]��"�֗�i��~���N����Ss��^�۾�M��0;P9e��D�J��A��`�
��m���qL�L"�6���6��z��c��L
�ea9D5��J�Dn�a��X�rB�D�|mj/J7(�/K��������zmh�������!�{)���O�]��ɕ��hp�l�
�+��PnK���'��!i�)��0�~�Y�6��:Z4`6+�\*�n*V��ZGtrV�_��3�6�E�'��"���t�48(.+��;��8��ϔ<� 9�J�"��Oɨ�u㜼p�=�i��ڕ�k�j���W'�	�k���#��k�ZNa,!����c��M��$�B�ہ�]"��A;A��٭No�-ۻ��@f�hz���?��H������#!i��2#�Q��V�����M;�D�19${wd9*eȾ
������y�8:e�|�R�Y�y����i�c܏D��tT����S'��:Nҗ��}3�Z�_6�$KB��G��kG$Ͼ�ܢ�i}���b�W�yr#���M�����2�P�gR���m�F�Э[W+�7DaGc��U^��M\9x5L� �������Y��lY('�qW*���YtY��3����)�/!Z'gU�`H_<���-�jAK� G��-;�7�ʳ���R��V5�]r�`�yl��e�L�5��/�3��#h�[�l,��L�4��f|ߨ�0���>]�Q����l����fጺ��gP��DVbV�%Op�iT��ȹ1�%L���w�UTK��Z��mÈ :�(��T'[��#{a��,�������t�W��̰�X:;�^�~���7���&��GVDLO�'���Aj�� ���`�"�8FFr�\o��	�����ˁ9��}����ؒ�Ė=�����%��VӨG��3|��[�Y��J5�4�}�[j.>�,Bh�ż��W-��:���ӱ�̂oh���喒6x�؆���˒Ը�e���k�4b�%p�ؒ>�pCEp�u�t�:���{{0���{�c�;O�;r��`�^R�oū��Ք9E�V��pX|�ҧ�PLU顉g�^�GeXܮ��8i��@�i�X}�_\�<���V��Ԋ��^������>"�nzz����ЭH߂�W�}��c.Y_�!�������7$Ma_z�X�X�:q�'�Q�\z;В� �D� (�5ߗT���R���c�����[T,���؞&��w.��&�Z���I}�U��	2A眾�q'��Ӈ���U��~��]�Ε�����ߺ�yNi�.d�A+�mnIぽΡ�4/���(�l5@+��#2�ެ�3��	���O��$z�n%�{�����z�c���<ps�+�~��!�?��� ���P�WB�������h쑂c�E�#�(��,k���#���˯�bNB�e�o���9����<�˦���.h#���q����e��-�U|�!?���:���W���}V��KW���\�_��G�dd������W��qj-��0�W�8>	�Cm	R�e�f�o(Q��Q��8�N+EɆ�Kg]B~���ϖ�%,���y}��Ig��ZC:���<�Ū���0A��Ù6�r/�R�UV�}�͠_O�3�,�,���E�f!�dϻjȣ�=�p/b��>�&���,dƼ��8t�^���t���vG�f�D���@^�Q� ���J/�5�tD�kj�ق��NѓEPg?S,"j���֫J����*(9x�b��~���P�`n��i_�>j8��y�Y�����l��2�@�s}rp��ȉ�c����B����ɘ� $��V�� ��m�}yf�#�R2e1`�%����'��]�,����4x���>}o���}9����.�#>�����'�Q�	����C/�M��[-�}ِ��u#^��X���Ѫ���V�7ص�	J��x��7��-��]�_.X���N�~ �4�`��3�����c:�6B)�N��PD�*p��B�׭~����J�J*�;e�R��F��W���^.���,A�b��V���g�{�ϸ�s�;krG���>ަ�����z;t����Ǽs��ѿ=T<��ţ����F���#���0I����2]o8��������Av@(���}8?��C}]����zy{c�<���[��'�)y���]z���e:T�Oa�UC��-��.��O���T�*\cGD���)b�)�Gȓ�@����-�ZnBw3^�M0���)|7�#,N��/߭���M= �w��-�0R��7���&���}!W'rg�W~)�#�op3��՝��V&ܦ/h*��+x��nw�<9h�p �S��9}����)�v��3W�{�����'7y�K���'mJ��Dy���!e���*��(���h�*�[��?�9�9ȹؠ�&� �^-�0������	�izn����]o_�H��n��!���=Z{H���yYP���A��R
|v!Y�h��x�?���Q/dv�{`���}I����.?��5� �����6U�hBr!#O�y�TQV��@o��kQ�9߁kRW��yv(2�x�9�I�#�|�S�]��Xd�*&:�lE�����#���
a�:¿�Ď�/���C��>,�]��4���r��Z�������l'zK�*m��բ��B�fm~raު=����.E��3�	.���n�o��5W'�I�`�J�v�8{?�/
)��P<�B��z�Y�\�_��F�P��R�!uYo��}]�>�RŪ�m )�Q�\"�M?z�L��#���V�YӴ�V9������v�ʲtI[N���m�E_�(|=�ڮ�3x�Q�P�����a��Τ$��A���<�U!"EC��-�	�����ԉP�Ǐ%��*<����h>�L6��;��?���X�n���~;w�~�����ܲ-�)_wtZ.DQY_����Ci1��j�cg��P~�^j��=)�Y~�`b����>W��@�Ղg�����_0ҸDlߌ"�CY�Ė�U�HJ
,����
�C��	`e�w�x:���Q@�D���z���q�q@&O#I�A\������
��Y�V~���)	U_^�
�{���7�'���f?��\{�[��z�梪��`�����Pma���Yp%�[�$�2��q�\#A�B��3����@@9."��������ܯ@B�q}��g�7�bJ����9}q�(�˭�/��h�o�z/���n5U��l���3�>���y���H^���Scf*��Zj�s����Uc�6:���u����[�G�����~��H��9�7�A��sz��5)�0�b����z��[$T,) �^�qW���jû�=e�(��A+�9N�jψ�����a<�� �6*~Ӊ�<������CK0��[Q}:믉�Gl�����rDXV�7ݛC]����l�m� $�}i<l�x�_��Z�d�q�ͪr�(�J�6�s��ǔ��p�\~S�����w:�u��X ���(�;>��9 �����>}����1��_�״ݴVm������C84�T2G�U=͋<����$����$��j�W��].q�Tp�|��N�:J��f��)i�7_�u�y��	��Hh�v'�0��8����'�VG�8I��L~�7��O�����X�cc�q��b�i���C�.�]��Y�&<�=��N�*�W��tn�$߬����>b�y�]�^R���rQ30t8'��s��W�1�l"PѺlz���ZT�H�.^l��}��y%~n�\A��ËLa�j �4�O��vn+��t�M�Ҵ���P팟o�ڥ�p`���̰xL~��̞�b���`�ˤ+Ľ#�"�S(IȪ̀L���}mp�M=�R>�eQ%7&E��!��|�	j���RW����������5Z�9y���k��?�1_^���_��X��F�A<r̓5�[b<�\�Ya�x�;xNq2H&���'��xU\W���{md�Gn(���A��y��r��8�ˮ�c�)�v��n^�DT �� 96�#���P��ݔ�E4(�S���[���a�%�����ֈ�m\�0�&�ڨ�[�y��!T@���=)�y;�	�RD�,��/L�������@o�Ŧ1���Nݡ�� 	���:����u����B�m�jL�'��~���:�?�7���cƢ���16s�M$�H�a��X,��ZSͭ�5��є��7-��HF�pE]d�xٶ���ON'�"İ~��=��jpa�o���]m���UD�}��}�6��ጫj��<JF=�ڈ��L6.������d�
��T2C(���}]�����u�{����3|O�5e�E�<�u�-�g��<�e8�����+Φ�C�%#䥚i��Eg�^W��au�c��N���TdH��z*����+��\�����np����mఌ!���*a�e7�h@
���N��
ں~�K@��aC6#E,-����E�:��O�:7E��P�7�|�]Y.�x�1��n���]��k��'~#�p����װ�-G��? ؐ�_��z��t[����`6$���RW��S쾦R�1K�� $��A���+Z��8��q��0���,���V5�t'�>'R�����	�cJ�`���9b�����g�?&��҃�*�PsN�xʙ<�Q�F��爠`hmd.@f��{䱍h~�"4����f Ab��fe3FMP"[:����笶�@�t�PF� 1B�����6vi�P�����VZ�^���΢�b\�5�@�e!��G(k�d)'��AM�߲y���deX﷘� �D�6��#�K�M//�	�||�C�N0pُ����,LS�>�e�w�ЎN:Oqq?<���[c��)�^:�b5�Y&�@!�s���GJ�x�Z����(걥% �.���=N��46�A�?�,u.�
�of)Q��v���Ov�m<��Ǻt7�#�:mFE*������-����v|�T�ӲlUqxD��pC~�\dT�U쏼�����_���!���V����9���3�W���Nk���3E��坹��~U�#�<��f�׊� ���>}ږ��z�q��ɶ&ܬQ ���f6e��<vڇ\&C3K�V��Jk��.Z�t���#�r�������;�>M�٭�`?�Fc[�������@J�Ux8���	W�.�A���w�%x*;���$@�҂.l���u$5�F������HJ�ط��ㆸ_�/r�N�kH�g�e�͊�Z�JZ�j��ns�j�®�дk�]�d����jc�aoA�
v=ИֹfL��v�W	\��*&RX��f*�G�]�7.W��M/��p�H�Z�Pϔͮڄ��A�u&H�VDٞ����#{�._���PTs
q��	�����j��R�u"Z֖T��B�wE����U3��\���s��U)�nM����WU�&�ʅ}�@oA�><)��6�_���}����{��2���*ޒ���]��;pA��#�񟎜[���$���ќH�?�|VBU�]hbx���?UX2�����#�j�D
q:�P�}��PM+�w�xnLSSO?��Z�Ĵ��7�(cٻd�?�Tz���k�ꨪe�l ���4���Q�P�7>XS��5Lʹwdѓ��8e��Ӯ�q-�
�toպt��%��=E"^7o@xZ��y�s�ͥBg\�8��q�l�L��S����y�V�i�`̷�X#���0PJG-��
*3�(����22���s����X S&����^�ǥr��8�2E����=h��u ;�[��m��ON�I����V�Y��l�{����9�D��T������,:����i��[.�|�VCYul�Q�Tt�?�-���E���j�N�B'��%0m�������2ԩ�����9�IH T<4���i�K��4঴��~�gt0���Z��b�,=����N�tdC)��L���`�j��'��3J��wN�,�Sk~1�}ϥ(od�r�}��੼�gG��Uqc�e'��0���G,ڈ�8������8+�'�!���~��]��i��A1S?���1�&ڗ@�Ȯ�	ٽ�nj�Y�j55d�e���#�5Ӱ}�����\����|���;���vƫ�i�lK5�M�|?���CSn�k��Lb�Ns��2����"Ս�9�+���){���S��g{�DI��3o�m��)���*���#qցjXҘ��)��z�/Ҫ-R��Y���ri�g/�2S�k�@�{��`F��{ ~��Js�1p(�&w�� ����d���H��D�T�z��9{ӡ��)A_{�H�n8��@��ɛ�o4@�����[s7�:X$��YH���D�B�����5�f�=Х��w]mY�U�����#ɦK�K�6�_W�f��10PG��I��Y#0�5S��w0�)�#RW�IǾ�=C�����6�h�s��&���-��?B���x���eN���Z�Q4|��.=W���G��y��7ɍ6$�@K,�O���q$ �} ����A6�G,�vF@Th�9P��@�o�#7���W��;��ꗴ;���l��y���}/4��3�c��>]�R=$n7T� ���@��n���L ��Gg�LW�L�Ӗ;�S��]BH�f�v�*�i�-ڦ�����*I��Z�v����HpCb�/&$���ѡ�;�P*�v��:�l�uD�J�	�Rִ���$�6xR�Vq7���\w�x{%|N��\�5y�]-��G�9����%uFx?�%�a g�p�݇�v'���r��E��`̍�ˤIt;�U���Q۝ѷC�E�6>�>)���y���zqo���I�Y�*E�2��XR���P��G�Y�M��J#�oz��b8v�N��5��3��� MN>�D�@1�dRh]ř@�6�����?5Z� c/�a���$<Q��Xx�iկm�B��I!SͿ�5�蹶�0�e�ɈLhmd�Rs�5��2��m8*�$v�rv���V��5`���З1o:C�]���y��}�z��y-�<�eX�뾋�M3��r�պ�ȋ1!�g��L��E?��yy�<a����4�3F�#X��i�P����hCFT�����[��uA�P�pZe!�IߘdX�����u����{���!����"�S\vx��#�uF��w@$�ެ�34�b!%�m�P�y��=��G�2�]�3�c!|E;ӈ=�&Ǭ��G��ٜ��𖘨��8�)�s�&�l|$C號�@�����hnȎӦ�@��>���K�� �hh��'�0(��k��^v�9}7W��z�uD�DF�J��{��@t�y�@��r�3����Hg��fW�� (�+5JT#��v$�Y�#�WB��e�ȸ ��ʩ�KKz޷Ѷ`����]�8�7������x�`������yBƜ���S}��>gK���J�dR��Nu��[�K�\R��Phο/� aX`<���S�sTx�q�E�)aٜ �����I�/0�*���mNs֗L��4��&M��uC�ݸ� ���]�O��\��B�! �;KT\<g�6s]|`�WG�#���(���|�ͥ~�,N9��V��wd�C�˼�ؖ�;�_qKϣ���)��RZP΁��x|�@��'S����/ >.쫉Ǒ�+!�6
4�i5N�����,�w�鿋荵S>ٮ���46�m�8$[��WWT`���O�nl����>�h�D�`($Q�ϱ ���Z>���+�Qܔ'�W�d��Z�9��T��˸_�d�`
��.�.�G�����>�� n=�NX�cI��������K=�^\(�����X9���b���Cʡc��\`;Cd��&���"�3�Uv��#f��$^D�#���S�M�lNt��e��%���qy����ȅܱ���������EϾb���O�0FE��NL1��.��P3Ɨ{ �~�s�M�\f�em�������-_����ѧe}Vg��,����I?z��	�k����њ�9�]�Z��Ob�{��O���\����%����^����/�4�߁�^��Jؗ!���f�6��Dt�o���h�oѮ�I��G�"�Z����+~��r~*}�u����,>�af�p^y�Um��-����kH!m�Gv`[[i$|N0�ڴr��ض1 ]��-��~�*庨�����V�����[y�Rdp
�.@�S����_@�BЦH/�v5D��χ6�1(�+�-QѱS��Gy�G:�	�RFH!%��=��{�����ph�A�wt���xxJ�)�Bw���`u_��u��B�����5��:SD����\�I�#p���Y3���Z'��ʴ.4K��e����2D1>O���$ɩLJF
qڕ���H�*�]�O��]��l����V�\>V�4�.}:1��cV!��
R9�s��(f1�`��ז����@)�����ïl�#�*À`�ƀA�y��ܛ��:)�T,��b�/��Cԅ������A��q�+ܘܩ�X=�"������*�gͼ����Фʝ67�0 ��P�خ���?��<�9�W�ھH�b�v�zW���xK{�4I�HHo%��ĸ�H8
��x)�L���NW�,��c�ɫ���9,��5��W����jU,�1¡����-���b�O�2,��W�?�!$��	�ӒB�q���d =�6·G���R��6}�����mm��I"�2|�,��S�*9�`�(S��sΣg��Y7������Z,�g���=B
^ytlL���0�&Z^�w-b��|Dz�2`톨t�}U���i�lIH�B��:I$���X��O�C1��@�;����&Gpa��K�f6w���� �}' Б�w�x��Z��2�"Pm%"�F������q�p��)��&��?4)��ߝZ�q��B�����zC�Q�h�q�\U�&���D��`�U�hKQP�;�6^����vhn3@שɐ�Nl?ͻ�7�_�����ӣ<5� �����	
����%�nY@�J��R ��^d ����'Q�P[��E��9J�d֡|XD t����`9��p���Mʎ�zQP����ޛfrɼ54��C��O��z�/S3w5(jͣ��p�(Ґ��;}{�.,5����5 ��>/O�����ފ6Gc#c]ȑ�R�����j� �HuVL$kF��:��䧿K�4#z�ӄ+�js̰M��h�8x%�Ya����q,gͤ���X!�qC���	ѱ^%cEb��6������.*[$��Tj�>>�DC|?��0�RY@ �#��ﮋ�#POSz�|�w��9y�Qbت�jb�X��O?c�R�O%�i���`P��پߕu9�IKK�
�m; �#���yْ�#}���<�1�ֳ�NC�-�0[tî؈
�����i_�M��> ��t�.�8XR���6���*�#��8\s��[��S|�,f,����f��6�p��d�v�je��<�0�y\��rt���I�$���Qitmkd��W�~E}~3�G�|ǜY��`�w���2��M����Mmj�}���7�.[K둊$�x�|B�됷f("��4)�~�j���G�~pA @��dY�sĕ��p�.�Hl���q�i֘y2@�����k�xW����Úb\�vM��r��/c1<m�|�=A��Q��n�*<�tXz�Tץ	��LQ��/m_�q�Ɖ�R<}��9�)���|}��ʤ�럤)t�K���������}%��[��?�"e�:��ez�Iq"��0x4"����N��h�������cF��Ϫ����ע��)@��� v<�����'=̐�NA4h���ʀ����hP��ǳ�9f��q�;��1=�����N~|�1�cA�"�rl��$!��|�k��.�+��X���d�-]��b&����>E8}�Kr�}7P�{+W}���SW���]�?��#mˌ����M�����)��D����r����h�t���i��I؟��=�{{>N;���2�9�Ԟu]��^P�������6�1�����P\'�+tЉ1��B�&�ĵ0r���zN�,�měg�o�Y�,�����ѻY��JSú�(bf�1����k��k���q��e��JI���`_y*x�cI�HW8��8I�
{���h�F��e�!'Vf0.��U�K����+��D��b�c[�o=���γ��H���oj��mH������$�s���l�5�{���9��i��x���˙�S�������� \��"ך<��Qf�W�}��0�J��-����/�a`��"����}��}sc���|����돟���  *��OX�+0��_���);�dhV8�С�љ��.�z�=�ȯ��J�^W��ʘɿ���W��r|sJ��e��ޢ��x�[�L뻬����式�5�6e�[hAF�vL D�r�[�����k��
�� [����T�$8���Q4d��Q��e8&����r�#Y{���bA'�mm�S�L�D<�#��Z��p�V�q��A~!ur�_�7�G�l��ʡ~7�C'��J�?���^�)E��DN���aϠ�n�ƈ�#j>^�$f�.t��9���5]��\����G�d+�v=�+�uݽ#S�N��h=�w��\���a��/��M��,���]q��m`1�ᚻ��~J�'���|�w��~qU�V�+9lт�zuS�ޘ�~'�٢uE$ �y�_��$VfoYO筤���2���=b��c�D��3K��R�opqJQ8F��Q��=�V�:����K�;�3�z��p/8������~<޹����ywl;�5:��G�C��5\��d��A�e!��ѴLւ��V��R��Iw?�a�p�#����:��!�?���^��9�_�dL�q���K��7A��p�bQJݐLiIF��eo�e���_��G�h�����@mS�^�Ϡ0��M����^�@��G�G���_�[s8�������<��弉�Xɴ$�Y�R9����;؜�tg
qޙ�CMȬ��I������R)�}��{m��o����P�IM.���mV���}K��ک=M^�@A9W�����d�l��@��k�m�&��OVΫV�_l� s���c����`'`ڜϖӂ��457��O�!�ߧ������W#��f�Ol���@_��$�~*oh:�˜�ѲH����ߪw��d0��;\��2M(����z�Xrid�P��Bz8�V��h�_XYoAf�^�Z7��\��bt�!э��Q�p��$��] �к��.jw�?���9K����U)� �}!v>'H��c׆F

�I�s�(h��S3X����^���;�m�P��\̤Y��>�3��w�̹��S��P�Ez��;Z'�p(�2�lO��Z��(V�fd5��Y���EFe�MxSm��B/��<ʀE?FHF�Orm� �I�N���ت �`���;�z�h�E_��l����<ۛ}!.ukSL6�;�!��h�C�e9;��\M{��g'��[�BE�'}D�z�7T<u΃
/��{�	gx�ؒn2;	'Y��*&����'yJ���iX\wO,�?�4x�jU��[B��Ԋ������pJ�?Zg9[c1&m��<�w�Nq��E�)-����!�T�e��#���l7f�����*q:/��>�T��X����K���}h�J9I�ꝿ�U��%1=���e�f�p�j,���`��;<�ˀ���8�K�L�cDr�_�(��}>��M=ZD�F����w�IxS����,�F!���^E
�����z��B;���������S�&�ߝ��<�u&�L[~������E���=�l� �m�,9�������O�h�闵�����ܽ�.1]�SGgj]ȝ��Le�Ht9��09�TTz>I��O�ʣ!kZ�!�GWf��H�<��:�I��a�
�<&�*�E�Qj�w��k l����b`��L�= @5�]�a���lUz���Q�ݷՆ���Fj��F�%��V��2?���kcˎ�Yt���#S��n��lB1�&%υ��Ϩ�L��aRe�נkhU$��};DR��t���P�zĶIͲM��1#Q0��~j�G��W"�+�Cll�p6V��'�����yO��Ŝ�^��F��å�9UQ"����v��z4m��/�_�x(��p�*��Wrg���*�����0���}�myPv<�Z�뿍cQ F&O�������vz��@��4���RA��z�^�23Lce�����8l�	�&��4�'�f����^Α[J��BT�j�0�]�H5�k0�S�V�JOE�#�v�M��d�d�%��U������W�+-q}�t5����j�z�T#V�F��a�G�� �bI�pZ��9����L�$��h�n�0`�^�eT/��=h�D�}#?��qI�|�'����E�f�V3�_N'rN��Ag�s���� I�3��le�\��:G�,���&��.>��r&1{m#ك��&␺�_�Cy14�Λ��CZ��X�R��V��ʑ5u��KKV� �g(�"T�K�u� �Y��Z��Jؿ�������9bo�N���r�I�`��ӗ��ܷ�Qd3����9w����d��ZB�,E��Z�}�:ٕaͲ�����+�ٯ�xAy�����:������T4�lA�%��IY�q�C����9er��T��/�0����#I�9r�5�e�6��d��-�T�M�޴�!�^ ;��yΙ�"T�T�>*��o����[O���@R[>��(��9�&N�"�����'OQ�����6��#�1s$�ҹOI�xI�:�9F>PK<չ6�r�^�Ѫ\ѓ{��o輹�5��y>9-}������ssc��۪�c8���XW_�� ��U��{���ǹb�O]����gM-�����]�`X Z�>X��ޅnW�i���R=�,4���� `o�V>���?=�����~�iLq4��)�l�W^�9��V}����*��`�^P�S�Y'���-�( b2�\��rKQ��؏�sm���B���Z܄!��'��)��X��D��bGH
��{n�3��˃�U�����cU�R�& t<�Ϭ�*"K���W*��_�n{<�����! �vXFHM�_�7v;av1����݆q��+������M�Y��c==�#|�Hm1��0�c:bѐ�� ��d�7H�d�_h5�\�A3���2�(1��=W�P�Z����d�T�[���,�g;�X{~�)}P����u���f��27��w}�/O�����_�G`'��<�F�#}��'�<e��Vꄈ?����E��6�]�5O`��nQ�>֫eŴ�-:�آ�St��h�U��y��ְ����<]��2qy`�ѹh${K����\��v��ؙԚ=����o|�saC�!���$R�{v�$Ml8^���:����-��N�r�(TS�J��@WRO~��,j"�	�\���w_�i<dd�ăNI�@ 
:��V�����FB���$�QQ~�Cs��� �(��s�� #��6���شjYP���-T*�z�
���w���	I�}[���ֵc�2_���Iw���dQN56����ޔ=)��z�gW�l~~2b/5
# h�{���x���
�, X�)�π��5 ���+�'�L�KD3��D��,_m���UD;ٙ��Ʊ�z@�g�P7E�s�,pZC¡����Bm�����4aR~����)���[�p�.����n9];}0Z��Z��\f�H��݌��؋��&~�s3�pV��/f��-�J�BN-k��+���iF�F��~����y�I�o��T�=���4�K��-R�c��pm�X��2ُ(����WH������l�zhb�V���W���7��H�8YV�ԯb�({i<��M���8c�s6�ރ&\W��9q틠V��v�D�֋�´����5w7�E�����A��30�Nm�i��TO/Ԝ�Y����,�Pl�&T�5�K�;�냙��и�Gt���<Uk"��G;���b�������|^$��C���Tއ�t�g�-�"ͅ�Hı���cO�.��~���I#���a7� ��8��~�#��MR6�o,�Y�FDH�N��=��o�6���z�:aE1��(i�:�,Q���U��$����t�d�F_웠��nrG�{yv��o�*�[}�Ǆ��(��g��I$>�&wgRό������@����Dv}/zm^����r���8���/�:��:�!��L��й{Ft��C�Ak�!s�$o/��ϐ����)���ۡ�b�xz�!a�o�g?���.=��e2R��� ���Z#j/�G��3O2	���؊�I�\�M����[�c4/�l7�ŏ�t��KI_6�^<nx�U�:��c���ܱo/ђ.m5�����Y�K��:�۴��d���5/Q�I�C�K�̲~� �a~�ɘ�1��@�h@X�)��c�e�՝�tB(8�;%��-���E��o8oPf��P��)J<���7��T�����f��������w�!���f����̩�Ԁ%vJj��iSd����w.����k�~0���ΕϚ8[S�K���v�/Q�y�/�Խ���Q:B�M�+G;�>Ʈ��.��.�#����]Ċy��+:��'�F����k��'Ut��&����Dޕ6yf����Ԙ}�H��f�Ч��}��ȱكO('z����J��?)�Q�׭̓��c�G)-Z���;���>������� iN�;������}��������a�ް
3Y̫q"1:s1�-�7��$��z@�䷔��^���ӟ�)���'?�	���Ӏ�&��Gu�KS��B�����nQ=��F��D��ejb��p���ElH�*W�<��j�{Bf��sy�SM�7*���V�������v�x[���sC���*r=`ǭ��$���Kq���O}|@[öC��vV�LQa�@�r���]�}���D��%���]�aI���	.3�����;��)k����`������>�5�����*�м�0��ŽA�J��&HK�[	�'&'���%���J�xbn�"���-X�i��wL���)U��X�?��ےdN�0�r?��XH����.h�d�jtq��J_��x]�1B8� ���� �����`a12�~����@B�r�m��p9�V%:���\���-��~��L+�4�S�Ԡy$��ە�P��ǳ�so�(�Χ��z�w����^�;�ؤK,��Y��� �p�t��r�����\����f�R���(��`#6�O(�m	ȓ�̑�	`��tL��,�Pꇣ�8Q}�3���s7`�P\�DVV�����Ռ�^ �)��kE�h����3Ԋ8{]�r�Q8&�D�P�gcM�8����ĝ��Q�%�\y�ZP����фC09?�wL�("t�fD�Joe�D�Cb ��r8��P��l�7��y��^�Tl��_��E��l��-��u�D��Z��*�����r�Ya��dg����ك�����[@M/�M���(BHD>�A"� ���)LԆ�x�+ba*%=���C8u\8���~���uC#\����۷\�zT�-&��D0VQ�V�e#p㖟Y::{�����U{n�t�eU�J�0�Z���q n/u���q0�&I�<~'�N{���VT�[G�1������ڲa	t_ߥ\�tSk3z�G�2�M"H#/���߻��@ؔ*�z�]b�+����,�Jc�I�Jt�thѴ%�n�z���4_�m����H|��ϭ����9^s�Ft���o�����v�O?�|� �H6����~q��q���2�n(���	��]5*�(�/i�����ȓm]����?���9�ܫfxd��G�I�L�8�R�jރ��	5�ߣ���}R�4��ۅȱ������$8=�*�.����ܑJ8r1�zf^r�io�q�e��b�@��"I	��^�yN"D:��k�'o0��N4���ϩx�FK|du�)�������4�{_T�I�1��MHV�u�N} }�,Sw���bPKEq$W�#��7��V�fI��+���QϋF�"�bwx������;k�=z}�1/Y�!�S䌨��٧h��Y�k�!��g޷C���G�s�v�K*&G��29�"�ڟ�)������"Ũ7��H�~���-�����z��#Ry�EC�l�����GS�l�bD`�Mq��5�߄쿕D�u��� b0�.�<���z�6��j�9�j��ޔ[��B �)b2�� ��m��$ݠ�=���!k޼��#�A�����''B+�	u��c�^��z<po8�wȢ<��l�9?�����j׈�k������f ��i���aL�j�BB�G�����\\Œ����ša-0ɯ�v�C#ts���*$�Z��,|�O��UoU����ɖ�?��q���)$��0�8ZOS�NqW��Y�,LM�;�$��0��n�L�%7������`#�	-��X�D���1%!b�̋�*��{z2i9�g�qc�0:�mm	������0 *1�Ot���<MCl���}�FJ6T��#۸H��X��&`�rH�M�D���]93��i��\�q���-ˮ����8S��G��2�Ӧ<5���ǥ�²�&zG��h 4��Bm8�V�g4��Y���&��AiL=��.��!���q��O!_���nE����U2hk���O^,���WN�F�%�T�C��^�S���;ɄL����h�J�K�tr@��.�9<�I����!~/�G���.@�v����e!���l4�O�������S�a�k�o4������g������=���8b�7��4QJWɲxc(װt���4�h`��AI>1���r�rB΀�57�V9��j���qAL�9�?pvB���I$�<b0��qN�{�hũ����H�Q�=���@�̯h���`2��$;�X?	�gA��8i�A�n���w!�,�ɷ>儧������%j�&QX��P�*�/�vvGir�ȇzТ�Ċ�`/�T�
�J���c9�h߻�ߨ�3!�p��+ [O��d����Г�hC[�*��˫`��ٜe%v���,4g7V�Q��~��z��#��".|`xe��rV�E�~꠮)�p��dc�XI+u����0q�ʱ��.)����/yERa�R��=)�ՠ��,=8GP�#��Dl�g�>:��n܊�� �6�j��d|6�#92=���aL}��3������S�m��ǃ��	E�:E�٣���Ҵ4�VZ���H(�SxO�Q�3���P)'��r���?e��h_�J/7����߷�uRݬ��E{]:=T�����hu�%*�V���l��}�$�n�Y�h��Eܑ�#z��L��Z�NW�����s�p��qGfD�ɔ�-l+���E�����qտ��7����� �]2�U7�D�T򜘇Z��\Og��K9���ɹ_�ؼNn��Y�"���֥q,�-(��L����<
z�h��W�����6�@SH�&����[�bM\�ˉ�Y3�����fYb�}!��0��%R.ĞF��.;5���F@�L_��!�M�W�j�dX�>�^�m����S��of2��S��Pμޥ��b")�0�u�<������>�q�ў󍂥�)����[���M�b�,����;���I7�h�]����Cg�j��2�u���sU1�!bY7�|+��bkZ1���`��rǄ�h혵�ǲ@��o��̽/r��VWv�h�ܼd+H}���g�u���V���<h�]@aW�=�~�}v�a��Q�f������Mpz%�ŬZf�����L h��ns�g��	��MP�꺵�R�=�]g*@�@����W�!�L����߿w�C7u �������E��U���N�R������Y#�X��]�-�g%Tn����7O�O�l�`�i��7? �L��Jk�0��.�$m�c��� �m9A�Ƕ=�APC���{�FT�EޒR�(M�q ��_|y� <;���p$�3S�R���v��wBu�O>5�e����Av[���r0V��~���;���!]?���v{����r�\�>ӈ&k;��尴�Z
2����
��R�����Y��䈆_�� �����*;����!���˦����b̳�x�-轎����榘v�����������{��s�?�>��V>�C�b^�A��cީ3t"��:�ŭs�vĈ]��Cќ�`ؤie�2�����ۚ����,�1"£�A��_ ��2���*K�Z�ǳ��*`h@̀q8�Cئ�S%P�'��*����<i�`��D8~ ��g�s,���[�Bw,~0��%�n�(�#���.��=�w��r͌��1ɑ�5}����:Q��8lj���^4�+zH�T ���237w�@�Q�%N�N�=��_�N��Ȣ�[�Ę�5�t��� ���� � Ѽ��͠79��_��4����y�3[�\g�U�7�(�u�꓊j Jd��)��$ �X�i�5�T��4,�h������'�<������aԩ��Ͷ�a50.ʕk}V�q|>��MWX���WY�*�=�]�	��q�,�Gb�b�����v:0>���@�XB�0��`B��UV%x�
V�[�X�=�%��1�Y���Fצ��y����p�\o�nC#��R�
` �2L^���}��Sy�Mh��-������q�2^{�e��,�G�d��돉��x�nDk�/4p�5�x��y_-'�*;�����p���9�����I���Z����]�IŞW�u1�Y�J~��ć��F�wj�����~%z���������lv�gQ֧95�ɅLxߋ�>��hw|ndxj �No��WN��#�	��fL���P��+W@!�O{_������N�}�$�m�1���
гn@�o2n�@12� �X���D0���+"�����n�?G��\υJ�����&�A�T��1K�c)�d,j��H��!nQ)!��#���6"��M��`�y��nH�aioFz��=��MJ޽���>��yb,v��Tr ��Xi�i��>Q�����Qt���;h����vB?�*���Աs�w"q�5��Ltv���╉��$J�`)�9��ވuH���l�}�)��k�S���D�
�_��1Q^.޳��;��}e!yU2��z����y� ��^ٕ/����=T�����m]��Zh8r��:������u�3u�r-�8�V}�ɭ�k�!��+�����@�~y8�''I�m��,��}�Mn��ടW�SZ�oJ�����#���aY�)|��y��� KC�{l;�|X\�ĈxS�p���B�����众�>
�s�w3*m�����Lp����;ә�t��J	��C��������(3�-�I)HB�����3Ħ�ЭLݭ��#���;Ӛ���Gn"ð��@� 2�<��J�����~��[����d9��!-�����C{�/Ⱦg����h��<�_�)����c�D��#�q�t����&�.Fr��)�&?��[�/bL�{%����˂^�����^)�)
���cѬV�z�و���Z�	�$<HDX��Ӯ��I���"��H�&�DJ�$���:��u���C�ES�U�M�8F��E�J���ٻǏ��c �������H���Et���%6��O�ye2��k]�u�'AwM�T�*?�6����/ߴ����J��W� ���9c����!����yJy�E�`n��H�C��ߥIɩ&i�s@ߖ�l?T1N��|�}�&6�Q������𧾔w+�{\k��ؒ�P��;���H����Y�j�ӫ}��cL��K�m����P����j���')��2C�k5ֶ���?�x�W�B`��V�8����ΐ݃��-yb��q��/9ūE=����3e�XMW���y7dgj�Z`��Z%�l�m�E�][�%�O�XK���Iz	u�,�_1���>+���#(���5C�ЛE>��v�K�E�ݮ��9���s��<�:��C���+}�����?�i&p?�g	�VǗj+�������b�C��t��eCǴ��vw��3�Lۖh�V�n_�>mݹ/��Y�h]��a��6�ۻA��R�i�rgH�+�'x��# EԤ�~�Ҧ���=��1��ܹ�m��ps-!���^h/'XV�Y��%��e����i�Nt���i�C��nw��"~a�b$�C�*�_N�MmNr�)���A�1�@=.S�a�&���",h��. ET߽t݂�z��� �z��[�.]���-51��8�A�t�Gfc40��J�BH.g�i�/\"j�L$��!����eX����Z�C#����h�Sޮ~�`�C�Hxdܡ�YNK:�*M>b�jԓ�r
�+GJ/H���ad��(n�E�Į'x�/�k��(�6,�j��d�cdVO�&�< cS�(�f?�_�S�T����r��
1�,�wN�����'��xWWf��h��]��9�3`*�+@B`j�v8��Nxт�򥭢[R9�j�ᚨ�HE�1#UݮnM^��6�}=�G]o�7������l!_�`eیP*�B�SPw��&a��Y�)��(M�Z��7�/�Wn���d��!�˂U율`�¡�#{%]X�C�#aJf�ɞ	����z�*ٿm�&�v�"�hfC�y�40���Ƕ��W,���0�#J�S�*Q��t%|t�2m��U��jjVz:��xhy��X��#5��������9Ch�7��7��"��:��'��1K%\L��	HX�mCĉF-M���Fm�ð�U�$��$B����<�)�����C���rX2�7'Ju^Q2�)O�1q�7�OUoe�� |t��{-N��o7��鸽q�01#-�;��O�\h�<:6G��������ޭ�m�<�WHJu��n�Jo#���Ǟ��
C�t�R�:�}��T�#I� ��u���{��5��<P΢��cO	��y3(���:�i�Dlb=^?ve.��U	;�/�ͻ��o�����j)�?:.��F�'ݝ��|U��p�}(�j�H�~�_�ֳW5c-�i8|��c�� (1rv�s��ͺ����t�/�4�?4�qvh�M�?����-����е�5�הp�ОF�F�@f��<������A<��Y�mPͲ��A��� �oK*�".ԇ��T�ؙ�ݪʮg�L��ؠ.���rq%��u�{���k��KO�{�CM�D̳�M�Y@��;.\ty��F��~N����t r�+��|�E_C�9��]}:�x�U?�H�)�Ҳ���-|�	�~�e��H�?�Y>n@: kgx�Lr��T��87[�$���F�|D:`w8\?/���-�*����5��ȗ��X�;���l���ϱR,B�}KBr�#�lͲ��q���#O�<���0��z���~)\�����N�V�������p~}"D:�a�����Ȝ�{���)�-��5����Pח=q��n-2�|����n���J�^��gXN�!�*F�+��p�L�@Jd�5"Ns�7	�~4𪯹��륯�A�s����& �b�Q�}�1���tS!���y׶k�3$2��Dr?�6�ő��r�e����ħ��P7	���F��+m����\��%������!��0��]�Y���U3�"1�8E{��Fxvl��7h�����5ֶ;'�&�"�v���i�	<GvR���#��ժ����?aK0ECeW�b��/]c7%�����u�ֲ�Gx��w��t.h]��V���YW�pY�iXAYJ�F���2J.5㊑�6�d�5�kU��"�@�)�����?��׮(�e�_����eGp��N��]�|jl������(�5Ug+��1'M��i�tg����ʚTK�SՔE	p��������y��eN����B��S.��$��������Z�j8}��!������"�Moas5$X�D���L[# �W3����W}f�2Z2�iD9�d�����G�?~T�yh'��xGoa�LĎ6�t���t�|R��7n��o�����8��XcV
����d�wd����TM�tl}-��|p�p>��l�m�+ɯ`0T��O�駫1�:��i:V�3P�O��e��