��/  h$�p�̦Rcس�4����&�r'���!�~�I9�$��|Ξ�ѕ�.�ߟ��#��&��C��u�y�B����=J�sbOEIwi���AXaE���F�y���F�j�9�J`�p�ϣ��(%ӧ7	<�6�|��Z��;�3�j:�&�㡐K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<��Q>�����.���P#=�a�3s%�J��B��TW܁�_��D9�`����q��?2n:���S(ݗ>��MW��ɶ�q	U��k-�p�C:ԐH8NL.�Д�Y�0�Te��bU Ln^�.>�eW]��mכ���k2%(�N3����C�d��<Ԫ&҅�\S]�k�@�U�t��I%�L/�A��]�L\��6��ۘ����q�����bSt�TԘPe��>❕������?Pke��4$���%Q�����6`�Lш=���/c�9R.�?u���;>�as!�;�Lױz�?�`Y�����ƺzNڣ�	���РV����V(B�� � =�k,���/�좵=�d���=�2�(Ҭ���L.P!?�wgt�N^~R�a��O��r�;�vj��(QGdO"�~�@�Y5Ծ1��̉C_��R5����"�f�&TTŭ�JL��^0u��e�&��U��
�FQ�>���Y#+�/�����١OܐQ�z��Bs�H�a�8�ޟUp�l���	g;=���&{h�!`�!������Dr(��k1��v�<�Bv���]"�}>���w�^����˱F���ܰ� �:M�>�����y�d���c���7� �����^E���!��
v���ٗ1��0~J,�1��~Y���a�D�XR;��8�A8�\@�eBu�}D�S��<�Y�U� �zb�&J���I�Fv�[����Si;�� �Kݡ\������eK;�N��a��2g�&�E[S����P�����h�����$6J�����y@�ː|
Fb^^]�`����b@>�����(������Wu>
�L����.b��?��5+��X���K��+���>���K��F�]f���rISVԙ�����<6�mb�� �V�c1&^� oR��kL৾�9��i�ja[I��|�044���j�Fi!�2��}���H��������u=
���� ���\HgS�,��O�7YL"%[_��G�u�Mu��A��2$ǆ��б��#����Y4��[ZI��959�.���_u��-6o(���T�!j�2�4�����xD�<��k
��,u��z���1���ے���Nx~ӌ�Bxy�֒<�륱�����/�{�O�*M��Z�Ǐ6F��P�b$�%�x���~��e�)b��D��=�I[-y>�GC,�(�z0�����`yPe�A�^oTQl�64A�\,����L���X�$/��[WD�u�s~��f�u�s��/��V�i{uA��a����2#w������J�W�\�^{�Y��C�Q3ava�:՛e��	vS�L$��lH�����y��b"a��v͓s�n��+�\��5��h�q<�[���1�O$������>?�ޫ��E=�<�n9�\pNB�g��.�ń\K���jk_� �,Za�۴�m>�ƪ#OG\<����[F�����B�8�mK����te���i6,������E��$�8���ɩݎ������׈n��p�40�λ`{��Y;0�ٔ�'N�aPQ�]3��Ҷ:���`���?�a5L�|��N�>G�=���xJ���:�{�K6k+;u|��㙗I6i�t�Ԙc�J��K+�� x���g�B�R��W�Z,_8�%z¸����?NK��Tȸ���-�Xq����/mxV�!;�l	��W��|��۴f�Sq�+�ǖB�����|��3gR���u)�zca��?t(8�lw
�}�,��{��4�������B�>�ϸse�ί��'pٷ��� ���Mr`��5H�Ί�'�k����N6+��qĴ4�������Q��'�Q<̤�������ޒ��0}��B�T��� \�EW��x0�b��y���� ʋ�j���V�������ֶ��J:���x�Q}���;N�j+c~iQݡU�|i�|<h�-�Diy#�Íd��g���8�5��N��IKӵ�v���B�I�y�8]b��H�=ӳ60	vD�Ogb��Jh��P2��Ly?��� "ʔ��V-�I�W(�P�Ɔ��ݵT�-iюO�6J�w�:�/hce@�vFl�1��ģIsԷ������s�|`���=���
uft�Z9�?CD��|�u��S7���b��'�8A<�v�=H�sd;�3$�����:���5/�]�> �ԱLER��u��ѕI��Vk���0����y|-*O޻w�%��3�&���1���� �{Bh)��3�|%���]A��>�vI��x"��3B��
�=5�+�x���>��ƕ����!�ׇb��[S;C�T�%U�lY����A�%��w�L
^D���PV<"��CQ��_K/|�^���Eu�C(��בl��8���y�HB+f��<�n���-d����,�#�~�ԓ�T�K��Bᕗ��fq�$ �5����_�9h��?�t�.�V�?��Q���u٢��ɪ�����J��&|"� �`K��m�е���Q��%��uUyr� �����1bd}:�UO�o���6~]�ѕ�F�e�'\��qY��X"p��X�0"��n��˅,[R9�2���G1�?�Μ��	H�=��YW��8�y���B(� L�*��6E^���,q��!���Q�SúZ}�6s/���d"y� �EAՈ��/2�y�a(7�__$,�\Y0��(���bs�K1��yXJ+�Gݛ<���M��7���X|\��e�~��'��dݭ����-���L�Z6s̩�����wʕ�+���eVH���oğ��Z�W#
z�0�=zV�ZԱ�߁QnǸS��,�"�Y*�J��}��LH�(P���<�W��<��/��،}>��m_��.�j��N���pȎ,$��W���p GO.�6�3uMR �	��H����a�g
�����B��?��F��$�������F,���i�,���j���n�!���Oy���5��?$ 4�%5*a�
V� ٮ�R&?�2l�DWt�+j~�H$�J矪Ka�u���Xj�
��G��N��|�pxh'�]�ϟ��I�D�%��EzV��������lq
Y�(e�۔����9���&�Z X6x�o��cD���K�����ˡ�h7#�C3E$0�]��KS�_#���	��"Z�K�P[,�g���@���?�9��G�UJ���N��K����AR5nڦzG~������x���I/:+�'����qo�o����+��읔�L�C-m@�ܨ\:;�����C�<o��Θ��5.�5/h*_���Qm�eL��۾c�iL�6d�A�4�������h`�.��l�jW;B�"�tM�l<�K��	^���IQ�ɞ�c��8�d���-#�@�_��CLm;�ډ���*[|��2{���b��71-��ſ���f�p��'�ɜyD39'H��'	G(���:��_�Ɣ��p.��|�~�w��XJ[�WE"��03>E�b5��	&%� =�A	u@��R�ILq*�������2����=�]�6_�u�Ua!���`�9�������~�����<�u7s8F߼�kH���N3v`z�'�ʩba�-��
���ݽ������q#��Y�I-D�a ���8�����3p�|�B�g/����W��
�-�	�9�\ۛ��@�����I�����o>�U��k`RS�zj���5�g=}N`d^�RSycIz�fr2�٣������	T�щ$�f=��f��/66;�������U�tۨ�Zz���%��9�WG���V�*�2Mm�n�贻=o�7�����]b�Ԟ��u�T/�Oܢӈ!�w���2��#L\��].3ˈ�{��K+=~z̅_�-)[�h������z��O�4�)j�v�k��ޞl�!l)����cu�gd�p)���ɻ�ٓ��M~͛࠵�l�����q�	�2CJ�̀#��%jƨB����Gb�+���.˥�e�@���Y���I�f'x���?�W��ll���ӳr��H��x���W����z8����~_ܩ�K-z�"�L���s�[�;.X�܃qQ�� �<NP�f�;��"+Q��/�^�K!��!�V3e��AM��T��3ȋdI�Q�~���܍;7��/�`/�;8g/BaK�m�Ա�2t��ef�� ���i��C�62�0u��`�,�s�,�i����+K'S�N�qt�<*e�Y{���ܺ�Yӡ�~Hl��+�;�E���*α��2�9�_�ǂt�7��z�؜f9�"Rp�NNT�;��Ib����_d ZH" �xsz}{X�b|����T�g�(e��?oO�h�[�K9����?d��\Q�B�S���BNxׯ�Sa�+r���RN�#$�R|��<��� �f�"_-^ZbO�,��lV0��k���D�t�:S�<&���ҽ�!7�n��GS�*P��DZ��]�*;@�K�pf*!�-bP�>�z]��Et"
��W�s�C�aג�F�f�_�*�<�4Zb�jNW���+��Q�lm�ch���,^:���Y��S�feC)T%ju��s���ٟ�g;�k��k䘆�ѳ�g|f&��h�i�~r��a�hT�28W��Vꤚ��-�х
`�.yKG��D }gB��n&���������P"��<��c�b�\�IDtK8e Hp����6�&�8���"m�a�5��໢���ݗ��@0/�s������ٲϫ��>��|���1���5@���1.�.w�F0ٙ�����D�>�����b��ٗ6��7S5�p�:��w@	�\�Tܑq��#��b#�y�|��OX�>�W�������琕Ya47��HFmOq9㎷���"N ����9��?��U: c(9��tu�8�H}[�M���..�ښ���z}�t�S��c�ZE�#qP����u��gw;��w14A$�p!����I����1�/	��k����P�@�r7 Kq8���K�m"����k	ξ���dwɿH��"��D�+-�f���F�%��GYD�k�޷u(2��cֆ��J\ܽ��c�����9;˻ʍ��A'��Fo�*���UF��\��XMT�����q�Hs�k�`?��w&V)��%h�~+g[��(�K(o������&Z��}mͶ_�Z.���G����G%�H"����(�u��o���u��̽:P� �QVI{�S{���%��tܳu�=�)IMC�NBH� T�-��1����R��ܘGؗ�=������Sa&��K��̻�nmNUO�/AMKǲ6"���`��ɀ;�F ��)�._�rS�0�p��»W���M@��6�1�LN��:����<=DE���ȼ�&��Z�N��uBg����E���fߡcWd����@�j�ꪲ5#."����,v��@^V��6�EH�1ʯ1\��`���]����jy+�U�(���L�K�BJ�w�`;���Ju��SK�* �ZB!�$�%۔�t.1�F:.��&�!g?�������lx΀M���HW�2o��f�e���ʠ{"Lw���-�$��É�R��6�vfm%3DI���.��{j6��\�̖� ��Fbq��f���׳��L=�a���"=���gRy�"A�����kϢ"�8�x�J���wܤ�jh���j%�]4��ȱ.�!H�J�Zg�$��J�����V֔d,�f	�'���vք�3jN�SUH�0�.phW�1��2I��qO�mʥF�_�W�<"J��L����)T���WCa]M�p��N��iX�uKXW�ө�߉��M�p"�O�J'��
�Lh��p�d���7�I��KHz�@�:.M��ɷ��C���?�����5]28�Sn㥦�6LG;2�$A$
�������u.xc��ӗ�Y_��`W;�!7��1F�V�J�O�z�#i�q��n-��H�?Zl7�G70��IA��x�:���(n ��z"ߏ�"���C�5�n	�P�ۢ��@Bg�e�y>�]�b���
�KRs�zRш��

�4�|r�����7d�5*����n)3K�Y$Lq�/g#�OY���kލ�@ͮ�9/b]�
$�յ�n[6_{N�g,�D�>_�ߜ��W2M� ن����R�ǘ�!�e�(0^��kKw��A*�\�1�M(����L?FBfS_���M_>����G�!d��}��iWrgRf0#��5��IU)�X�U�r���R�S�h:o���,`�i(���栻�#�EL���x�:��!�4�~E
W;�^�Wq&�j�Uza
�b�&F%aw���#��ֽ_���?��0�8�X�{}l1��RO��j�TH�=��{'��M>�簼3<+N�h���V=:)�|o/�5NQ۶�p�-�Ka�ckfe�6�N��d�B�3�5"���?䪗� �+1q*J�z �7��n��ù&+-'����x���;H�٩*�{�ݠ]��Å,?���G�H��DL��wb� q?�|��Ѿ��Ҙ��	.�M�!����]Ɂ&f������E5�Tf��%O)�K�}[u�?��9Ԓt���y��nn�C���}F��m籘������' <�G��>�k�����t�?��s�>�aSʎ���(f�vm���0!�v�1e��`,��i?¡�e�(_K}�7�:G���T��u�7-���r��Qa���e"� 
�3�d���dd�2����6�"��Hne|�Ƹ��LL��#��g����-Dؿz$��E���(��L����g�EeZ�x�(�`�ާ�Y�m��١>�ʲ�@�:5܁k<(�0�x�J�v���W⸶ً�ZP�5C�P�q?zD��>�����Pq����%�N�d�L�Q�8k���q�8qxb�
W����\�f�z�n��h�4:C��]��=���X� "s�i��܁���GM�h$�\��j�3m:�W�����p��:l1�����,h�	"����$��U:����j����.x9��>��ݞ���pg$�5�)�)��AG��C�g�Ɛȶї}V	ŘJ�?$���-�B�0�ô��iX���s�2����L�=�\qԹ�3C����)������5=�L)�6����C٭Q�(=i���Q;A1��ϧ�6] ����m4$�b��X�']�����ӂ�ݝي�$�=]���3�>NMnAn�C&�P��ܥ(%�])��_��p�io�b^?A�J�Nf����O�;��<�(��$�xBQ�U��^ ��&jb�|�X?��?�:�z�Ѳ�[Q8�����|��P|�k���C��<�$�߄�	�{(CL[�5(�9~l�5�ʞ{�HK�*��[�T0?��?U#�Ԓ�U%�U���(��a����/�L�0���Fo,n��6+�|�РV�(D�,����O��q�u��ql��nF+��\N��K��,Y���".���و��A����"-��ڢ���;�ũ�`���c�`U'��O�H&�|��u���x�P&��|~d鮋�P�8[g�͋J�/����W?4�p\�̾��
<���m�E��AzR�J�Pm��0;au�0���W{((����[3����yG%�h�8&v�Z����$�P��LUUwc��s��I�P�h�5a{��{��M�X��bB!���n �r�&�K��,o�B�f�.�k����>(��\u'�7�נ�\[����W|O{���:i� z��/B�pZ}��A�`�27G`�3�M]gĚ�U�vbl�#%I[�=�L�e\
M��"��KPu[����x�Z�����G���@�ɖ�d�EH��N�J]���l�5{ޖ+��pA���d��j[�$���V!L�Gӗ9��IJ�o���r�[C0���~�`U�r�Źr)�o���w��!��'��
Wq�c\L�J��V�(�lۀ)��è��-+.E�J���v���>̢+�����u�L�v��xhg�}�F3T�(꤂��=��~�iw��[�Lo�d�˝ J6����	~o��1�9�;ΝE`K�{VV��/�]�-�7>+m�bВ�[%�_����?[�$�����K��;$���ŭW+��o~�n�8M#����S�`���&�~��`K�WcIS;s�aI^��025sқsƟ���[����[���7���okh�M+�	�Wd]�Ov�r]��۬51/?w�E���u�ON͗��ىK��ɂҼ�F׶9�x��DGz[e/�ґ�x��(�#�i��k��xR�۾K���=��^UD��vQ]+�O[�~�]KFOc�j@S��_p73�K�C�*���6:B�gO��iƩo���7�wє�B�h&���!��p�P�Q�_��mIln�$j�{ �j�%����/�Y�N�f�g�c�t�x��b �Ȉ��o��.�QY���ar��qC^vD��6ie�8�y�,D�z�
��&�ߙ���g�87��*<Pc�� 8qY�*�к��])�tZ��t�lo,V�)�-_�s�( 9+�
������B����.�$��=h�J������G�%n���r���Akh2[�(��/�XT$ŧLiJ)��D��M}�а������޶A��d|\�k��� 38��>����L'*z�j���[�>�N��ʲe/�j�,.*�����F8��O
B)!D욤s����P-0��9��IF��D�5Z	���⦂o2}Sע/�VJU��k����d��H����1Y���\J�N=���Nw�w�B
I������qG���E�X.�����;{��2�C��:��0Ime�b��+��ڴOFJ������1�B	J��kB��os���?���� w�)��'eA��+�D*�̶4��j�^㘄 �,
�1�N4�G�]���;2VC�΢s�E
(&��)�Ѥ�!r92p�W��[!�\n�3VHK�a^ݵ���bn���h���W�O�Bt]�}$���mQaX�ɥ�r��F����������H��a�2����?.�QN�h������:/=K�2)�|b���~�`��Н���5}��~�v�X*q�yr����40Ţi�@�Ӥd �.>�~�V�Qs\�7�d�w�=j�rչ�L�C�`����H{����s7��ޓ��b�;����r�P��n�)[�{,��/���}��Ȕ�x@�y�|u�Û��n��m?(j"�O���@��)�2)�㬻w͛��_�|�p�jǣXd{����Z�8�ᕝI�Y��m�rǊ�)e�w��;����$v1.��X����#�py$�W��)cP:�M�`V%����$�<L߼,���4,���6�b�A�/#�