��/  ���#���"0D�������^��P,������@��u<��<���CQ�#�����ͩ!�]����{>e�z��T0��v-|eE��\�/�J.yw�Al^�|���J�On-��
]3!����~姐_���Fj�,X�T�H��!���L�� N����18��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!����ıL	���dG׉:�v�&7^ș��+�W1���_� ��Paj�u5�����Q��ߝN!(F��2!5hv��/��1���=�O��]"��Ǿ�Z�������VZ�����P�����;Q�����5UV|�`"�j�O����]r5[}�^;] |a��5Ɉ�x@���i�}h��̬M���6[f�ׅ�H@��f�$L��i�4}����O�as{`YJ���Wx���!Ǿx'�q��u�a��������̨�)��/��e����㐭���>Ȩ1^��fR�W��bQ�� d����[JѪ���<�Ӵ �tV������^��^�:���-�q��Y����4�l�d��\��>�Md!+��,'��]Ed� ��L���Y��Ӂ'��.���+�Մ�6����6� dtSA�Z����Ȫ��	g�&a�6��ܮ����	"��}�!��-�ȑ*O?A�B�L��6�K�B��2-������wr'9��w\|e�����tW"X��jT��:ij�a,�o'�el�+�"{tC���2�"����ɀ��#2��Qtc��\m�H�X�Q�Bܤjԃ��/�+{s=GQ�P���H��Jta��$��bh�^�G�}3|��6�
2�K ��YP_�D�5�⣭�Zر��2{#A������̟֮�5YO�̉�k��T]���LV�U��hz�2�u��o�/I$1_���Y�k�_��ض�I�֦�ܥ����f?f����,�g"�1��d./l�4ӭ�PK4�X���"ȩ�^�,��s!��y����@�>ۆ���Sz��iW[��YP�x_�0q8�������>��ӆ����	�����f�(D5��\�"N��;�B֞������F��s6��@s�\x��;�Sx�\���|*����u!�>�$K��S�	����A��3?��8|�q/Y��n�f{��g�8T~��Oy[*�҇W�q���'�ȟ<܀�<b��@��/�J�Ľbғ�0��EoP�-�9�s!&�*f�;��0{>Oȋ�֨�s�&�y;��6�ȯ��Ȝv�kK!��1�b�V�>,�x�:�>i��x�@��@�gUN��g��������'@%����F�nq���e�ؓ,������/	��~fw8uHh�J�F-�a��$���P+=�IÏ)4�1�� �����u��zpְ�KR{mn�3�ŊI��.T��y�@R&M���?w��Ѽ�*x�"������?v��7�Ǡjs >�l���K�p���oA؞<o��s��=�?%tJ��=)<&�n��Z+�p�������̜X��X�K�pU���l�ez�*[*���]�K8��L��ȧ�-Ѳ�菎z����P�J���+����
+K���Tn�)�
x�v'K��j|���b#<��nႲt`A��k��iP�\压����#�;?zKk��O��h÷�'�8�v��H��,U�v�7��Ba�ASY�~ô?��@U���1���H#�U��,�Z�dj��u�a�LT�۬�aX�26�����Ex�%Ś�����_ G�hXRS"��b�O�)%�{���V��Mk�q�e������+s�U1�o���>_8Žנ�����7�������;�R}�j�w%4<���3�Z]Cn�崈'I�6I�Өa��ۓ��A*���d�l*�3��A��u�*����aө0�H��cҩ�13@K�s)����ۦ\3��T�>
��sx�1�>l�'^*�٫x�W�&sךg�Gm��NA��8�{P-v��)����9��G��٥��ɱ�~�x?1W�E %��H"N�x�{�f�"=/��K�=�्�
��E�k;��ˣ,���XLFZ,"��D�u^�Z�c�U�vF��2H�`�\h��Fp�ߦ�J���Q�$h)��i��g��kAbu�&F^���h����������D������h�{H�{�X��� 4C���aI����T�;�Jۏ'a���*�����By�=T�j��2��F=-I=��*���}|}k���j�E~��A��u6,ۂ���+���qB�,c	o{���|�,��+�N��ӽ�-WᰓN�$QcZ2�f��01�D۟�C�f;V�0V��r6�}��$�� w��;E���O���6P'<��Ϡ7��$G	�{�����w�/2��;�Nމ4
ً7� ���������>�WGN|X�lw>�Q^���x��!�zz��tN'��@f3�M���?`�3zvs�Dd��=��o�!�A��`�F+�C�fD'g;�n�h@�X��0��r�:Si���?M�G�wO"U��.g������6y��ׁD��y|�t
�ϴ�'aN���bS�X�)�R��C��ڽSl�Nǋ�v��'[���d{e� ���1��M$t�r��;A��(��r�z�Q	h�@��4���j{^�ȍ��$e��a8�tL�.�Fx���v���nЛ����#�\�9�������*�h!�U-U?�u��'����^k���4c�B��LƢ�VF�s�iMs?�CQ{�:_��,�a�_��u�R���K�Hî�7�n��./_R�8-%'�c,�KuS.��8?��/�;�'���{��ޱ�N���+t_d�Cp>�r7�/=��ɼ]�m���@ZÑ��M��nq`�ܬPK����i��Uq�t�:s�櫔�ړ��fU� ˡ}<H��H��3Z���8-�����p_9�̺�s��
[n��g�x�c٧��������	ɬQ}����wֶ{.!|WGݔP�������ŨVCLb?m- ����,�SY)q/�B�5���/�ɠ}�y�[�x)ly?�L!����i�Fb��/{~SU�z2���#�.if�����Ao�b�����?��q�퇔��N!!��vom
�v(I�<��|Uj��
����#"č��3I �S�KW{�}���h)>1|�nٴ������g/�2$g�G#�27#{�$���b)RE����	a�c���E�-�L�=�Jr&��b��Ƌ�J���"�]����4s
`Lx|֔CW�ϵx=ZN���\y�3�K%S��L���5~��r5fu�<�0?��hZXmh�w����6��\M\�l�Ӿ�u}�˙��D:����o߬���#��G�� �Y<��&��x�������oU�Z����AX�`��XM���%>�Ғ��t�!�4ug���0��!�F�@g%/AZW���zJ�d��3ц�D4���!���#�B����4� ��Dz�n�q�����2�nY�"�����'rƄ~n@��~u���:�6	�#g�߭���*�ʱ�b�	�h��e�hV�YM��S�
K�!�i!D�幈��py
eo0��P����b�w�9U���������^xF����R-���x S:�k����L���_� �˓��g�fO����t{b�L�$Mi|LOC�1s'"cq�� �:|n}')W�n?f������`L��������F��^_�=]l�+���<�����ݪ�w:qo��x+�+n��:NŊ�տ2��O{5���a�"��$%Fl��B�4�&�_v�����^������Dy�k�����m��>�kUV�-?�q��]�ˣ<���3���3HZ��{��c������dF#,��L#.��tanc�c���"���c���H}�@o��(��sM��!n��R�����#eI ��o9:2���QF~@l&�8��������c������]LfTuE4(�W�����Q�H���I}���̹�A]�TS���a��&M뺏�^Qf�[C)���o?����@v	��q�IdH�0/h����r���G��r���i�4&��H�Ģ�N�W�Udy��'����>��{uMbK>p����W