��/  �L�fB��;�+�]s�_��&�DF�XF�3(59�\���8BV��ѩ*���}u�Ua�����)	}>G��Et�6SR/������W�.�|�D<f@�q�;	C�3Y���/�pӧ���Hv{�I҉���pf�>1�C22m�z��g��ɦ�ڥt'7��/^��<�J���6�����֕������h��3�"3g�Ĭ;�:.���ga�eAݏ��3	e��� �H���E;�@k�����D���83U�n;h���Xɾ�����A�xo΢{("�� �j��KO)7��
)�R�>g�L�I!~y��� ���妨0������AϤ��F�M		�?Ҹ����\��aN��1ŕ^�#(ƶ�M��=y���L���C8+���j^��ys� ��0z>U��t�\�Qt���S�7ю�e��9n�u� ���&���I$	����z"��8�Vh�G&�`�����d�v�|��tI����҂�VOJ�p�<]���t��v�^�!�\�Kw^�H�����fŔRۘ��f���W����4�T�(�M�7�Pۼ�g�N�B�ˁ����J�,j����������6��p�Z����o�Wv���N6����I�\��u��ix5�5Mİx;q�Jc�8n���p����,P <���� A��շX�t7�����Y�S����Q_���@�o.�%B˟{`���(H#��x���		CZ��q�խB���km���E�����9\�K�����ݒL[W
�C.^)����^�H�Uy�*b�!v��t���\�F�� 2���8p��r�.wH�ޱ<�d7�/
�`G�Pɦ��y02*m�y� ��2�6>dE�SUVj�,r:}�=t�B�<�΢�a-�'?" J�K'�<f�M~��x:-��ʤ�٩�b�'�I���bs�$X����	h��F��_�2�� 5}Z$�髲��EoBI���H�e�M��;���U���:���B/y,���{*��w�����Y��Y-������
տQ�i��N6��z�q����?D���t���re��/o~�>)n����q�\ĞΏ��Ŀv-�BIH'+;��Ը��Dn3X��	�S"��mV[1 ,�G�;^dM`�3�8:6��R���S�@�/���� ����Q�rہ�uv`�͚-&��ɢ�2��R�E���ዥ{a�����8p�W5	��B)�����U�_�á�7�P#��c70���y8�{���Bv~5 '�+q��&�%���� I~j�(ܥQ�`of��o�i����8��\�"+�*�G��XV�]�G�@	G)d�~W9(H������J��O�&'O1m6�H���e��i���\x"���ǅ]s9�����0W$���W��_U<E��T{��a��=J�@���!K=C�rE���Vfw�3o;F��P��$T���K����>ڀ�L�Z�L��zţ�ߌB�,_!$��AF�1Д�Q"'��B%n_���;|��_0���{��Hs"�e�a� 1���Q��'���Ίxw0ý&4t�2�V��D�5��Sؖ���DťMk�$�1u�c���!��77�c̓�����s^�X�c~gw�o������̧�#���ޥʵ�*ؑP4H<%���y�����kE
vu~;����F�:}�4� }�|&�%�j�N��� C�{.�u���'�*և}��w�K�D*�}��9]3@�!�e��+1lA���.	<@A0��{6������x?��Pd��Zc{��Xk� +�?�@(���ytB����������C���LD3+UN4���J�X�;���%&��̮/ �A��v� ��j�!0|!�!��bUB$-��c�#f��ه�)oVg�J;�b�y��Ƌ�xİ-s�U��:]gA5Q�/��_���y���Pr�֊)�Ϋ�<l&߃���:|��7��)��HV%/�3%zX�v^�ܗg9��>�k��!:�V{��@WV��>027�^�B5�ί�����eA"3
0�����:���޺� 2�����l�v~�r��~�<�\�����w��Q�V�6�h�W��=�<r�t�V��צ@���C${���]X���6s�n#��7q�ީệ�Y��xꝻA^%�e�q�y�aȱEC[9�%g
�r'�c��a��	�YK@fl?���m�؎.0���?x�N�@�v�ʠvUh4 !·Y_p*�����Ϛ�ֈ���5��OcVQ��9�����Զ��Gpa)�˻@��b���K���w8�ʌ?a�+�y�܁���<1����=��K���څl���U�}��ƼXD�eB��sX�t[J�՛!a�4��h��	�G�?�M�E��GD9��d�T�E)J?�`��� �9�X�!�sp7�E��W���)/�� ���BM�������'� �#Y��Ǒ8�F\�w��h�r~K���e�$+`@�nF��ק�5L�)���:�� �a�f}������g?��,�(�l���U/�XA�!x���b%?R� ]����et�W�D�B
��3Q6&b !s���`�� ��1�ȥt�zӲ�Q�Ը�>�&�R�\p��3��������k�	�Y��X��U�Ww�qS樚R*�#,�>S�se3�}�]��_�U�x�Qe����D[�g��][b�m=c.�W<w��-^~��b8}rB�����M�=����h�BV���֐���=�y:c����D>#Fh�ק̒߳�,�D�Ry�'C�8�gȞ`a:����SF��� �P@2dOQ	7���9�Ϡѳ��}��,`֖^��3Ň�����:uc��yީD�蠾��vt�y���3��DQ
�$���ޟ��J���\[�뼵{s�����5<݌P�yj����= �y8X����������W�S�,�֑���b�=���C٭P�>�!��.����=O#mf�ꟽ��!�d9��}��< ���j�aV�Y�_[!�M�L�Ҝ|T��w���a7�<H2��\ַ�?'Ն����V	�r���=+�0��m\|�&8��oPx���Lb�=D�'��e��n��R~�@��Ǐ�Qt	#aݹ�J4��ǳr$�����S���Q���1`��$�	d��0�質����(��,��ߎ���$��$	�K�pȍy(���k`z`d�k�n掿M�'�9��4�w��!l]|1L���]�r�Գ<z4�z�)h�:���	V�d�H0���]%OB�������`����`QI��oS{$�����5v��ܸ���r��A���#u ���)Zn�m٩����TH?��w?a��%&�dr� ��9��` :0��|�X���#���o皣fI�ߺ���G���s����0=a�p�R���-F<�(�T/�����@�O��a6� � %�(y�Ӥ��*/�#�O������C�Bt4��<68�ʼ �ziʍ���l��ݠuu��u�ò<�X��[�o�ust��&ވфy���P�╇��T��l��V�Oݙ�k����<������P���=��^q���������uj�fr3���^�u<��nec
6@~K�G��Le�@�����H����|�El��>u��-�hyL���3�r7��|'�Q���.�w����~�9��\ړ_�Ù��j�I0S�'L��n���ܰ�yO�W=���%VV'.x-ы��)�B�j&�x	1^~�\yAǅD�� ��)�ʩw}�ٜŁ����pU�5�b2Dw3 3��؎2�:�oX����k3