��/   I�����3Y�z��g�؟J�jg����a����b���̗4�5�B>Ȃ�׊�,��u#��G�|�g�T��!��:ۦ�ā7�"|xVYvG��M�0	`�u\a�*����Lb1�b� ����'�p��t��H��ʿ�/XȼWH���ژV�`��]ԣ��B�Ra��?rz�Ҝ���n4��Us$IBE.dL�0>��Ѐ@�\
��:ppզ{ 6o�br��Ҷu�:���9��Ԁ,v�W��cA�5E	����� ��Ӈ��8�7A	���ԏ�Q� s�α����5�:���'H��9�FfQa�^,o�g�C���Աl�# �lG�wE����P���q�����b�\OTv<��^�Z킔(�<t9.�+�|��Y��y���$�X<_Ȱg$	|j$"�<��<%+oRП�6�i��u�r�:��#h�|�������8��i=�<x���;#������>���XtO@\4��C\�#� �D�����GIo�dp��yq�д]=E�	����Rn�&b�K˰,-�����Vȹ�����a���]���)�8OP��N^Y��gs��:b������f��cL���^Ħ��A͟�������i�L���g�Q4��g��4�,����Ŋ u��کe<>����Q�"��
"�C�D)���[���}���n}��V[z���_�T��W��͐K�B�
�%��I$�M��VQ�8!|1t�4�������Qu�\�^w�4���ƛA��@�.�6d$"�,*�&#^���,�������J�íc�;��I>��	/���i�E[�O�=���<ݓ�s���8@������:C��PW�]]wU&��ybjL������=:K|7����q[K�-̷,���jy����~܍���Z:3X��Y"���$�$�`��%7-���-~�:"QiaD�c˂k�p�ڣ��y�S�����jw'g����X�<��Py��er
	F���s��4��{a�[C�n�PH��X ��s Q�]��2.����=��]D�T�b���P�w�SW��2L��W���d5	ؤ� )�q׿+u�"��_�U�j�eC���d��8Z���H�����[����t�-o�pe)k{k����f+�����_�#N����e����.������ͼƧ��`��@��˟~M*�瘓���}�R�d��¬�cM=ݾP�dI5�������E�z;���V �|u��3'�7Ðmw��L!���l�o�����
�\�_�ehݩ��B���A�W����7�����p>KXb��u��:�/��R����=e�l
�Bc�me=�v�y�<q+�,�I��3 ��N
���0��y�fp���+�^U�m���~��������r^#��>Mta�.&S��qE;�h]��M�P��ểy�;I��҅��^Ŋ/Z��KL�����>��_�2��؏��k����r"��e��Eg�<TVC����Ki987��;G�22�nT$�@�'W)�fb:t�+���-��%H׭��g�]��xDÊ3�߽�!/@<����;�qO�e��P���uB�fB���Y�uX��龜�ljr��z>wmnw\(�׈"��eD�%.%d�c�IZ�m�����7�]ho�����,�.������D��#��r
���UӫQy�D��W�dh4�r��s���7?Q��,tU��.rYvk��(����' �7���P�t�I������\��t+�m����(�L��~�<k�����&�!4��o�Ue��Ep�ڭ4��61%�v_ⴠ���7�(��A�X)8 R�WjP3�-�t��=��G|�dx�bH+ � 7�M�"}��������ӧ�EI�Am�N����I�(�2�M,ƛ�q'9d�����M�=���000�bR�?�x|uoY����k5!��U�����ăݩ�����>�+,ky_g�4���*!�Y�5̀Я��Q�=F�F�<o���
���@o�X*�'V�=���d�mT|h�y��
5��>�X'WP�+]�"g^G�A!@������]��.�;yӆYG�փ`.���6	�鈄�C��������s�{���b挬\p"q{�e_t"��"l̪w1C�������S觔7vhS��nE�"_�����#f��z=��L'o����z4�f��.�q�=��L��%�����;7�g���x�}ʡm=.tZ|��R�æ�f����X�O���Z����Bb�;q�����V�{��� �"�!J��#yO�K~��4��Y{V	������c�D#4K�I���,aZi�Z!S7�e69�\|r`��6o��V�U��&E��*�?|��q(�"����T7��a[=�j!�����I/igq?A�jKi�n#A0|��8���WfAa���g��|�ͺ��m�'9�?�a���j7"eRQ�ӏ�Q$�8+M�݈�j�:(�?�¼Q�jzt47�3��~ƾ4N�	{��:Hf���YP�|��:���-�LJE,�����e�ӻHs0	�;�s;��n�%��uFW�9��R�&�m�պ�����I�>�����p���.�S�BL4����[0(�;�B'�-�Kd6l�:��ͪ���еCi,� �gb#�~��#VN��`C��g���/rUȦ�q�4�%�چ��z7���a#�c�˦Q�h���޳�6?���O�IeD�i�'��3I�mK��lo5Bpث��dt'n���?�p���2���l������I����Fm��R:ιq\O�����`���g��N�g`j�� lS�RQ��jR�eMl�7�FTz�s�k�I���[��X���iw^J�d�VM� I�?�V�'�w9C��a�+��R:(��Ӑ������J,��� ���l�7MSE�cbO�n�9�0 X܀WhX��ߏtƅk�>I|+hQ��e��K�ǀ�?ߌ�Ѯm`z�ř�kQ)�O�������Q�"��)�M�UfxS  �͵��Dx��Q��� �`�^d��R��F{Y�,���t �bvq��|�ol�� �E_Ŝϛ�L-u��a�Z����|o��e$�;X�[���ӟ3g���g"}x�@���X�ʂ�7\&�A�N����&�>9��w�#4���P�4�r%�G֫�<ÄzU��� �-������6���F��t�2�V{�kȤ�;{�����U�˳T���X��abބ��HxH`�=�U��9����a�?��f#��|��ֹ~�߂��PeV���|�u�n�5FyH|f�����3i�9io��-�����{�^@vРt&�Ls\h�.D�|Ԯh�#��!�%/,�S!;�:�K��r8�I�%�B!�%$P�h����ֺ��66H��Ý�k��]�E�o���m��҆��&?��/ \^��_���c�w{�D�'h�=|zW���{�r������ޞ�`�燕}���ҏ� ̐. ���x�i�XT3*"Q��ګ��/����/.������D��`DJ��]�LW�w�A�����ܓ>���ݤ}��UER�;q���sDO��R�%l{�N��� :cPO!��K�5dR��/�ѩy�g�/$Ϣ�H�t0���@4?N�II�������,G��n��k���0��j�����i?�>�U�Ql�-ĺ��P�!)գ.E��9��Ă��h��g\�s�81U� eE?N$��P�Z���3��1�r�P���Isښ�����4��%y�����0:���H"�f�~(7ؠ�����=��Rӣ��a��0�b��_O�Qn3�_��,+�@;J(;��q��/K�&z����Ī�,Бl������)��;�d����0p�
�V K
�O����D��;1(�p�9\�wi<�8$�|)���/?Rp��*>��/�j�q�5�����"bc>���Z��	lJ���L��g$�0fl�ɐ5��]������3���%�K��%���8��V��)WQMAy����d��رk�dPg��{5lP���`�^�� a��>&�\��`/�����!r�1bWQJ����ZQ�iט&Ѹ�5���4����%��0=���9�����?�����XL��^��!g��
}Cy'�	�
�{��ܢ��xX��MOŏG�Z��-��0:d�}>�2���-+M}�A�%O0A�ν�'ħ�tt�g��VQL��j�k��=l�
�(��J�8yT���jJ��`n�a���J��L����He�ox ��YpN0<�����~Ht�cjʑ���Wo���6���9#����'�!ّ�*�ހp=.]J�����ђ�	-���iˢ���@��i!��x���h�E���Z��A/uF�3���D��P��7�U�+iA�hK����M�i�|ӡ��E�\C�-2Za��`V���lq�/gu�� ������ȵ
�f*��Pe�FS!�r��F�O�|��SS��i(L��H���30iC��JX��z޽+Qd��	@>��Ή������ �p����-�R|���x�B���A�nmt)C���	�+�[�e+���H` �b�`<�V��m�6����"�Qg?���&v�pp'(s���?;>P�%DK��TG$�7�����{m��%2i���.�{9��׶zn�mq;�����QI϶�|����oǡ��	-�>ް�K���b�X�nSd�w�WG�v[�#6��̸�âo'0v܏6�I�I���ˣ�ߟ��Cy��r�;F�X�4�9����X��^b�H�[zW[pGY��j�����sd�ֆVP�-��ON��z�5�P��������@XSz�<*U.��F�7�Mz�-�k�f���.���~�����ڡ*�''�S1Vj�����zM��z
W˓r�����~�W�ͬy�;�_"Qm��k6u�Tc��
Bg밧O�5��ihg�K�׶�g��w#&9�z���m�-��Ű�:�gx-Q����Xrl4���W�Q��D��m?��w
46�!��ǒ���ַ�"
w�ԧ8�
���ɉ��G���'�^�1�����	ƒM��)��u����NhB
��2H��BObF���"�Z����5A9�h�ߩ��m�ɷq��l��$�ZNA�D�AѼ���y�sz ��ŶA���ᷕlM� {v���eӚAƓ�Ԙ'����6��N� �07=�����&�WYYޮ�9�,��@��џ࠻��pG4��ҙM��f"�����2�HW��8ث7��ҵ م<�,^��CPA\�W�R�6��q?SNs]�%��]g�աWr%|��)��8� 2)5�?T.j��o�e�����{3�5�鿼��hHR]f=����'�.	�'������cQ��Lc�T��׃i���ӂ���66� o~��WF����ݷ�*��y܀�g�|�m�����+ԑ�֢<�~��������KL�7���U[�q�T{�Z>,���bH�"�+��DT'���m��ȿTU��a�9h� �R/dts��1h�X�=P�*Z�s�B��#���*8~�]rf��^;�73Q����fR�pM���P��!o�ɟ�����
y�L�Y{Rd˾a0�(��?�ץ�m�l�&,�mhv��O*'����Ҽ�l��D��g�7W��G���Q�"��K8w5$>Z�y�1d˲��}
�6�����n�����C���^"�_υ)mT�c޿�nc��3�e;����߄=��WO5�U&�x.-� ��?1K2#��y��b����!�=k2�r{�_<3]j��]���p�{(�_s����; ]a*ɽLBL���������+b��;��p��$�]!�"�IA��=�ߊ� O�H�05T����'T�CI&�5��S l&�_���-���!�o�{'!��v`B��qq�ϙ��p����u���E��$]c�D��.FWIb>*��R�2�ì.�I���%i@*�j�w2��@xr�߰,\M��UL��?Q�ȗ��9@�a�i��7��T+ae���7gT�+Ğ�����巬"�/�8Y6#葵�,��uO5�\H�V8���i[��aI�7u�2{a7���N�h|�]�!��"��I�Ʉn�O���HIv�d�� �"�/B��U<�7��p�^�A	�:.��u��S+3�˞���	Ă�f;ub.{;h
�a۲��;��m�^!�ϧ�ը�]�D��(l�յ����
�-�y��8�ZI����	!��h�EOQF¸�X�<K0�C�#'�T���Z����=��o�we�Z�|w�j��XJ=�s�!v�ɩ���@v������iF��?�f�}�{�꜅�J��Hx�[V��9p٭�	v�'(�:�J;I:�Y5!�����|�.�F�����	2���3�[!���]=���X�������ؘ`Md�A�Pw��L�aQ�n�]����Ƒ��ޥb�+
��Q�
�.�˴�b��E�ӵ$���B _ *�4�����>j�/RV�|F������^&��U2�߾nP��,I$�񸖹��m1�%ݘ�Xil%O)j#Ľ�����w���u]=�L'3\�����%3����h�y_=��L|7H�ԙ~�I�7$a�\��SF_*丯M�����?Qy�J�r��7�	�]�l�.�Y��W�r�}톽�<�9_��ߟ5�N�0��8KH�$�i8��4�}��|��'�Y�=
������S�wU��xJ����:�#��IJ�CP�0���[U��!�=:��8$KG����h(����M����f�.�������}�p�S��hC���;EԄ�D��
�п${���fuɼpIZ
�ş��ث|6�l��� �;�(H�Q�(>%�Eh.j@G�v��
1Pތ�V�l"�3�b¹W�]��� �<�f�6!��d�lMT�z�'r4�@�-��Ô!��A13?�AZ�b�7"�}��f׻$+����4[�%]ʅ��}�PWE�SrHBO���-Z^}��_W�R���S��S��;-������D�}��"���o�b-�K�w$�d��\}�Z�u[��Jywֱ�<L�^P�x�4��Y�(�V��g�����ٮy��Ҷ�2��T��t�3pzk	&��s��b�:$?7��pޑ�Td�%�%'ݖ�)s���&��% �.���4�r����i9��λhxV4��g[�"���Ɨ���6�c�X���y6����\��AfO�4��	~�I��=��6�pQ�{B�~hhj��p*8�Q�9L�eD���M��?����$�\+D�2��0B��o�ϒ�o;�'��q���^`w��#�`��awK��:��V�������ύ�g�B}�'*�e�~�ʟ��,	=׍�#dvnRn�$#xXA���ɲ�Im�G,?��K�j5,�W���'C���S�Oo�2��<鮚cj��JZ_�����1�'�O��8͟�0��,���z����C�Lb.�y-�;净�*p,�<�fd��)7�_����0M(��/?�:��Y���!-f0؝��Y7��6�mH���\{�Ne��S+$��g�od>�:e���l��}�?�s��+ºȡ/��$�g=�l��m����8��)<���{��{�L�Γޟ�h�t��X��ﻔe'~�C%���T�nۛ�4Y���5%}��,f�NUSG:Ʋ��j�
3S��+�Y�:S���������(������SU��Q��f�Q��58�꣚Zț�	�?�xo��?Sep��6�(�� ��k�8��E�reš���k�#���t���\\/�=Y�S�6���9�ј�?B��_%�T�H�4�	T��xإ	�p��������Y'5��J[�5v`�ɛWA�&�K��.fp��7���TJ �������m�+D��%�`N�Ň�*[�#'��1En��L��^�ݰ$B�`��qUYy�q��]nk����9 ی�8����^�g$��շ9+���?��Yz�֊?���My����̟/�Gt�,�>&�&li@�&������OddH���{bP�PK���'�b���^��A��X��j��B\�j���cH1.����K�5W���ga$�C��a�Q�\3���2�g�����
����_�q'�-��c��̊5uٲ���� .�[ʜ�0Q�ї5������b�N?��A�e����SA��δ�h�MIO�b�1��k���okO]�<J۴2�=��z<��W��.M�^�ج�0r�`�o/��A����N�2�]��P-R��K X����1'�^�R�[�n�=|櫲���cVc��&i�!�S(6�.�2��t7�����3`��>��Vcn���VUф�鬚�;��+���[�jV�qTS�^�k�����ttP�僫�`�sSq��	ZH��P���T�(�(��`<�
*d\�,F�b=��<P�ϧ�iD�C<m/�}ZlZJ<C�禅q�P��ː�8�D�Ks/+�T, U&:�XKʐ/ b�~~�\�F�a*�5��*x�Y�H�I��8�#�a*�_���%���3��<�TT������o��?��\�ɓppy��Gq�?Ҧ��y?���cJ��g�+5�g9~�䒇c�Q�L!*^�����,Kɽ=��� ����f+J+�u���h.
�9�U��m��]���;��ٖY�Hc)*A�JS����@�C�6��@kvW S/q&����x:��9cn0��E��J�\�3��7h�@tS\�7q���wu�x=�f�R��\^��8·)8@��e�c�RL1����7/�F�(��) ��Dl�5zf�w}&������^�$3\��2�X8@b�T��Q�sn=>�B����8dVC!��k��ng�b����|a>G;�Y��p�l�^T����׶�U�RZM\~|�̱�g��\q:�c���+.4,ȧ����������D�u�nsu�	5�h�B�S�s:���PA�ʏ�N�/�]�,y����r��c���Vt|�% �(5Y��D'��t����j^���֞�1�F�e���l��9o� �]J#x��p��ޙa)y�4_�Z��vqa}�g�ڂ����$ۊް*ۼmbgvď�<qmB�'î��'�@J���lb5Au�Ƃ��g5��W���'�f�`͢'�l>���C�;?��X_��~��>O�W�f�5��T�'��@��HsML��߿Ѿ���3�L�J�h�Y8��4��?=bU1�"�4Li�4��-ʾ:>��F��A��@�ϹhTѻ\Z��r�#�{�ǤgvmE#���U>�u��p�Fwvv����vP������䠲VS��팁gkQ����ϳ�҅9{X)�GBFB:���ym(Q32%窴�9�tف��`����Ƒ%�&<�j�?��5A:p���7���8�C$Dq��
�-�^>�u2�� {�ą�yU$������$Q�Kx����XsE�i����R=�`���Z$���A�R�1E!V�ʊ�qs����&�5w}�Si�&���ɘ3���Jܞ��52��c���� ,و2g�.�DicЎ�s�����#�7��Z�|��J0ځ���e9���g�u��{�],@)'!X��h/�H�h$oA/@LնAE��2`����L0%נ�F'�v~�Iȯ�YeU%��Ҹ��2K�T�6y�ٽ���Do�n��l'�k��e���+��h"!Q��X*�8|ߍ�B
��`/� �X߻�@��c��N�lw��돞�8̍���9�z[�ttO!�����jt��7ˌ�xC��u69�O/�M���4>�����Q�=�8*ȑp�J��HZ�VZ̦}�����3 :���>������6�Kj0W)T����A��o�����5��A��L�����(�a����t.��k�A2d���ŃMu��=��x�Gf��}:�Hb�r� "���G0�|W�������z�����B_U�`�7�����o��m2��i���f��j'�[�����iU�8<�y��������Ӌ��൱�n��ό��LME�_cP,��8o���V��@-�ȋ�g��#��Vl��`��{��M�5g]�Ə�8- �\���=�U�wE�A��3���z%��+ꇝ\�MWi�^"_��z���n�	?����t��K�V��lzhЃ��>=:݊�@5G��_��H�ƴ��X0�r9�u����Vd�54���1<�E��`>�Fb��̺�S��}Eʿ��F�?}�M���3���DTt��_�!� �Y� ��r�?��UE�$d�-�����\i
�m�Mk}��2|�C�5uX�8@b�x��7H��.KE�D���i�\���W�r�T��\9�k��]-	m?Mf�$�Հ�-1����8X�N�/|����;�!H��{Y��'�SӚ*��x���P7�3����JB���;��]1X���
�~�Z���k�(��E��#!:�H�uq/�R���#ڂ�YH_���J?`�� z��ڀa
x7�k�����B�l�Z|�����!�����T0ckZ@�L�i<�x�~:������@�(�t��;�Vb�q�\\\�ه:+^�^��y?�٫*�w��G�$`yw@	Tű��$����3���p����P�_e��4na(I4['lauo�IS�	F�E�tO��U�Ԁ�m���,"��	��#�rI�ކ��D[�b���-�i��fI5b��P6�A��N	����R��>(�OH�X��9>�N��3�		S�S6�-}-)����~��2���pv�F�*��Ŋ'����IH�A�0�'����Iw��b'VZhQ�ުx��&�'�O�k��T����qU�`�H�0DztV�W�lL�D��&���iӴ���=j�q���j+�IŌ}�gM��t����ԡnJa�J����g�Z��_��I��*�׹��hz��ۉ�m�^߿���,� ��Å
�Yj�g]U�9��'���������5e���<Nq������)���4|�-)�Q(�:����9�;�|&�^6���4�0��b
)?}�7�:
��U��%kn�e{�k��T����]s��@�=w�!�K��W���E�6ֿ9~�|{�Q�����GwYp�O�4�q�X��<��������̌�%$D�eEU���ct��B��3��Bm����q����{� ;�Z���='��fs)X��kYm��Gyu��Y9\s��Z�H�?�gM����j���0��QoY��M#��$��P(���ޜ��mˆ����y�����.���q+x0��W�?���4�IY�����}�Em' ��S����*@x�큲�/�H[�H�^�yC�Զ��v����866(&#u���[g�ؐB�ZF����Z 彸���H����ˈ�̖��,���#�l�P��i��wF�9s
3�h������!,a`�Fvt(���{d��� ֝K��:|�s��Nr��,ve�_��+�hL׼Eg#T�{`�4%��q=�f��EW� �b4�뚖�Y�ł�9�%�����i�S�e�H���	��\
�e%�&rY��X���젟{r(L��B3�v�$iѿ!���=����� 6�8��0}�|�z��ؽ�ާ����h�2e~Ȩ2�~g����mH<9RT�
�h�q�N�S]y2�����O�&m@`�Y*v6�<��������}����"��!N�d	�+�L�����ՈE�Dn)h)����]�v��p��:%r���{�ƴ����n?�D�/�|g�^6d=�bB�	��������F�~��0�P٪N���I�r�.�ϗ$KYܟW�V�ˆ�_l��n,��������*���D�
��ۈQ�?f���h��C� �?��p�G����'9?���r�f{#W4l�;����BbA̶� ^t�\���h�aa�k�{k��&�~z!Mk�xFZ�Ruou�n��Q)f��fî!B&�Lq}Q��UN(�9���� ��[u�ϲ�_5E|S~�Bc��8�����:�Y���3,W;D5�S4����U�?皪O�G��u;Z����Y�S�_��JCUT��j�5�r�&�v�X3c���i�˂#m1
ֹ��Es�J�,��o~#*�C�HߦC���d�$נ�\T�)N�@>Nl^�{��gI�a�\���\�ګ��Ȁ ;����P��m��P�ỵ�;�����%ܟ�PD��jJ���Q^�yC�Ry�'��x�]�st�E-�l�|�!�F�&4�������	�Ƕ�fݼ�ZZZ���{H[XU�|iDNد��{/1�}�|��1�SC)��#�9�bk���{n�}:*~�&������w`�B�NЃ9�ҭǜ��nsY+�_2��-�=xg�C���p|;�0}>Y'tJ��hQb2h���@�U�TU�pc޵�m�$���Cl*x���7�>�f��^VX�ɏՖo���
����3��j�uvtߕH�C�X<�]h���oS�Ѱ��3�J�q-_f�h�� f,��	��wd�r�b��X?���vx�t�W�P�ĩ/
|K��k��	���b�(�5tp=��6�Bkg��]S���Y{j�oy��i�2�I�O51.�h4�l��8"M�dFE������µuK�����ȓ��N��Y�����/W�؏5��L���?&��>����H&���ԑ�XPA�$Nڣ��7.����J��
�2Bċ<�����a��7�Q�l"�����~_jƘot\��*����ė�*�<��GC ��gt/��l���px�ϵ;D��#Z�w@t�_��)&l���<b�UZ�@�uʃ�-�r��=���ָ���-�������Q�v��P��V�׍n �[�s�Mu�uA��M���QN=�K���hQ���v�6Y�Rfq-�(�������g[4꽐	8�$���9��9�\v`gL�@'q��,c�d`s�!�ުF"
U�}�x���U1��~���aY�M�K��۾���hڃ�<��?ӉL8d}��T6E���)�]���䅪/�� ���&n{���i� ܪ���Ч>Ǚ�ϮA���;�7�����9�6!m&�|lĻ��J�Y������ m�dr��&9f�jp_��ɛl��f^fIf�*���A�����-��I����������
mOSo��7�t�n��^֒fL?^3����:���PJ0����L�X��~�|Yu�ʪݕԍ���w|T��`�T��T��]-��?�L�`0p�b=v����-]����<M�&`����uy6�cd#E'B�NI,`f��f�EKt� ����{/�������x��{Z,�j���mL<x���������nLe(��+���֜���l�#\���V@�@S�	0�PE	T�H��P��#�vSL8�}��p��U�9�R��*x��x^�!�ZI�]a��Z��{�e����˟։�"P(����7)pj��D��Njߤ���X;�J� k����PQ�-��O��oVkh�.T��)���"?x^Ia�Cc�U܅����2�>�F�*���C�'�q�mU�$E���X�Ճ�~�;���z��OM8�@^c�9^����s���W�p����m��0��@�Zv=�a�H���ۺO*�m��2��v�/��&;�����lpC^l$��5����fu�j��OF�ـ{��F��g�60�s-�L"I4\����aA}wOk!9�A ��&"�R��O+b���"^8!�GcRզ"?��q	�wAb[�tT�H��5�u�`����7���X�K����y�(�����V��;�%GE'��c183�cx���R���q����@F�A�z�,�V�8H�Q1�l:���n6�ɨf�Ё�PF��O
�B�2�mwF����'H��*F����9>�ݢ��~�$`)i��hRC�/��1�?�iq����n�n�����	��:+bRC�ʡ��X�R��S)�6U��J6fK�	��%e�Y-�P�j��M*�V�ۘ���y\fٴ]�0Ydy�S� gj�@H�p�?`��T�lj�����1��������cLS�9��� � ���:oE�pUN�E��1
�!�B�E���g�*Nvl�y	�
2^>%t5�5���UF��'�~u�V"ym��]e��"z���� #� {ݍ�&j"�Ø�����u���d�1 ����I^�l�ğ�좻UX�ÿ8^�� y��1�zE|"6w��;�G�HS������Asl���=�dP>=��&�T��7�s�ں�(���a������<>D6���f�b*3��u���7���l��� Vӹ͍�����V����R�l/���j��Ă>U�������9�=\�( ���4h�K:��3�4��j,l���yAC0�� l�͔mM�o�w�x�������=J%%��g��Xύ���2-��Ta$�c����Ţ�>
�N�|�e��U��6��˫c�4�����9����,��G6����V�����f0J�|�<W����8SyTVǰ#����e��c��\+m��/�~?s�(�I���I�)g���@S7�us������TF�nqw�e":b�zc�kW׺�����E
l�sW�t��-a�<���Ӳ�yB�����k�,R�"=�bjni�?��Z�^�PQ��v0?�ja@=�拲p���r�G�G�0�.a;�X%"��[
���or�\tM����_oP�r1�<Ka����#���H'����o:�\,�a
U\ܐ��[�z(B�^����¨/��|�4[�JD�7ܱ̋W�[���a]��]Ss��ɔ�4�;![R���e�`g�-�#��Y�ڞ�f�YH)��2�H±!rih�R����9�:Jv��`L�r�~#��ӧ�*3���Z���a�TY�	UUH�0�|��·2�r�yP�\�P����_D�� ��^���E�����t��~��Q#l_�G�큕�h��a�(ϙ�+�O������}�מ*Bu|����}��B�0e#��5�"1�����J�y����&��}S�c�	�>��ύ�N�D14ɹ�jvP �Lb����L~��j���t#Rb��(�&C��0��d�e�3;��O@-��>�c�r����a*jLPr�M��*��Cφ�d"���%R�ۿ#ҋyMnFUE)���5�aL;���,�ɓٽ��);�4��=NzL���1��|��l��r�j�*Ghue�v1�|��=��u>�'��v�/�[6P�����+�>�;y]r�0qr�R�R�̆C�
�Sv�i�[��}��g��O�#��w�zd|,��5�E�~p:�ߚS<�L��1`�{���O�Y�4��1�l�?��m�G� H�g����˂>�z�WS���>��̔}��)L���w$����A�:$��������"�7ϕ�b��D� c��� �ynY'�J�������y���q�%8Z�L��
��/�mS�W[�&��F`�:�)l�-5�� �E��xɼ�C�kLLB�*H�\Ȧ���dG6��L;��2��#}���͒ve,�L�R�3q�����2�_^��
�yfmr��Eg����g¶������y̍�@��Y���e~���k�l��j�
�O*���]��t���l��5Z�-aq��L�`#�^\p�R)�x=��==d8-l�R\�u�
q�����y]�{��%�?���G�ŏ�b���3 �O��6��&��%��P��lB��	����ț�~�7��������E�Vͧ��?C�çO�kx�������A$�YS�:[���T�٫�8o��J��pT�[".+��Qr�s��O�.Bb�1^��7��Ś�3<���x�+\i���]g����R���<�Y�G��4UXz�PP�n2He�	*��zgn P0%�κ�2X���&�*�붩׷�l��%_`Yv�yP?/�Wn����A
���*��hPF�E�������P^��Zе�/�-U�v���]���?�p��p��l�*/)vr&��k���O�;�J"��}��������م��kVc�c���LJ��X�`�qS\�4{�i;�vrw�6 ���]y*���z�0r+<��:.j�+�{�W=����?a�8�Ȥ�U0[�s=�22�ˑ״���W	zL����g���	h�������IA6�g���]8��D�#�Co.o�G�D���������u�c�4餏���z���R��(��+ϸ�6Y��TҰD	�	5K�y���X���q~}�L�E�]̷��Z�Alm����� �aA�\�P��v�2_����n%>1�A��0ə��"껤m��0�U����k�fHg���n��
�"%a��Vy�-��s��j��'\��U���;�I�=�t���r��i��z�(<�$A	̜Kh���]+ߋU�T~\��2y���;{�I�g�q�q�$�֪�h���(}�����ڠ�����zӚZ�>|[�>���S���pql��߆E��cI����?e�+^eލ=�5:�h�s>�Z^LU|x��lL��D%kE�ڔ������q�b�Jؾ1\E��5B��-�u�6��9u��ɟ�zv��ŘH{�:��Bֵ́	�*�'�ϿT�M��SX`��z�	���_|Ը�%�8��)�����ZD=���"@����{�v�V���v�z�������]�t'��>�����=I+`�Kw4ש�Xz*�7O��-7��7B���>� �4�-K[��� �blre����2q=�����KZ��d�wP�Ǩ��O����\�1Q��$^���i��P�Q���ƙ��Ľ��=�0�p�v��3y~̖>[+�n$�c�������r��I~��3��"�\{oW\�S���.�[x�"H�f�>K� ���6���}��y���ɸ��`^0M�.��m҆����֟�:0h� +�Q����9�Z���G��F��Z�9�3FL�5=�]h�y�����9�.x��Ě���"ח�}tx0�4�e���;k���	�-\�2CR`�g�s�5���7N1�j!�FS��)=�RX�Uic��Ÿqv�O֡�>u�&Vr���[TV�>1+r鱆0�]�����B���Ȯ �\nT���+�#���~�![ m����%������p�Mv�
B��X��8_��h�qIg��D��W#I���Z{�1I��-�Vu��{�'pw��l���`�t�kƸ��e�j!�C��"��
�9�����{�E8A1��x����d8n�!��l�D���Q��3����;��e[`p�)2�Rii/�xh�o��0��"�8�WjL@qy9<ʨ`OM"4�W���#�����S����	�ٖ���~�oHs�"�P�>��6zcV\��j�ſU;0�F���75��19��9�I�t�,6+�ۓ���&x1G ��fK\&(>���-�G��(�Ǚf9E�<g]h<��Y��G�h����G3S!r{������.��>p�c�Eˠ9Vܸ/���]#<���e6��}���U�3�vJ�j3�w/��<���R�[�%����6ԁ�9�Af�K���j��(5���@��c��7��Ď�G�n4�TE� d����jV��s/vM�����M3\;�2�m���D�S�� �]6	�j\��К��ڱXX$\��*�t����>�P3����g�I�]`Hm:��֏���bߗS��%(.�y�=!��Max/q�S�]�����R)]>��j�B��mK�}lT$��Zl�n�$-A�ݭg|�%�f&�Z?���C�`��=U��Ժ��(�P��
��3�F^��$}����)P��ة�N)���!C4��RZ5��c��5�&��{���@Ҥ�>��6;����PZQ�`����=Q��;�"��5��\%�ATE�U����Ӭ�[dT}x�C���F82��3�sv�Ei#D�E`�ns>~cְ9�Ysˀ@|^0	�j�MJ[�16r�ՇF���[Yb�1�98�Ȟ⧊t�o�""]T6�a�&���=���dr�X��Oe����ǲk��ۍ�R$<Dt�y�:�{�uuNF'�CXZ�]�7���+�gɲ$8�4�'�H[��ip1�9��H����7R`��4��=�����P�3���aZ��ϗ�nv��70�:O�U����z�����:�`�)~l\�nN�n{�o�d:^E�'R4������'F���n�6��e���y2WM1��<,�Z����I��e �i9��v����,
��6ƝR�|�+�4����n��r�,FSQ4e����íEv��/�8R��Lp�0e�7�|F�>�nϽ�xG�l9��읦`��(.�F+|)Nȴ�B�6�8���fq
<�&eѤ�������J}�ҔVg������
ՃYBv���늊>U�瀹@�N�6��4�(b;���9#��u���s�'�8�Z0#��u拯��L��Z+�MRbs�'��wo�Ig��Q��{��5{����q�z��LkW��Е� ,."2͠dG�}�Usޤ������F�'�����=8�[�*Pe��ҫ3��ev�-�@~Y�gX�H�4_"�R�����'t�E�������|��ⶍ$d-$=id��b�ʃ�P��V�n\ߤl�Rʂ
��t��m}��R��7U9�h����I�/�0v�q�*�(ȃ����&�)E����`��}�PN�V9J�]��Y'�EU���S[���NА;{6������-�8�G�jC/��=�|�~:�e#lI�1e�c�.}���C��{p��|�m�2����h�#���6c��At+�!�#���M7b��"j��b0K�}mף}�<��B�)���1��)!�h��F�$��.�菱mk�/9�[n��PE�P���D�j��/��(�$)T�;�&V�A�y�N�֟�����\�LG R��,����2�F0�5�
0\�k�BTaem�6���ku�G������'�!�4q���@W��qnU�$�mH��i��'�b	�����MC?�\y�0��J��xn�@���Y��?�F��=��s%}UX�5���E���F�GU��[��9I�8���ѿC0�P9�Uwʤ,Βպ��;�f�4ïw�R0��ãZbc�������W$*��Z���pW֢'��) r���F#��w/56-63b�&=k�$�~̊���&�D�]ҏ�3�H�|)�M)]�b]��+