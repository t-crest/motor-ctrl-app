��/  ��u��?[	�ȧi:_� ����GI.��]���p;� B���{�����I;F\��+6�1��H�~����"��曨��l��2�S��ܛ�&�i�*2�����A
lGʝe�Q��v�6�U��m�4H,�CeS �Y�]��w3&g�huOo�|�>h�
�^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK �7��N�NHtp�
��~�ae}��x1WrU��,-��ۧ�F�K4;z���� �`���0�N��<�7��{�4V������Yq^h�2�A�5��΍|\�O�Kް���0j��_O�s׿�XJ�E�T�=U�c`}�ʸT��P(�\�ԧU���z`�϶��~��re��Cl�?s��B{�܉|09�!�����8yE3�%�P[����"�]�����Wb��!�	N.\����=�w8�����U�t�=2�
���\m�P�����;;*�`�B�@��c��-�QmG������CS��%5 Y1�/Y��X(�pa f�C����S>�4�����D�l�!�2S�:�jA�?����=�à��%��5��ҋ0�
���'�@v#�o㰒�Tzv���ף`MV��<nR�w �u|\-��HY��K��2�%�U1�o�Ҁu�d���6 s�DE����:I�9,��6��:�ie�#J;&�v���)�!��(�a�:ę������	;<��7�c��h}����>��1<_y�F�	�����+|�%E�h,ޒ�a����Db��y���9|��(H)n���lU뒁�mo)�$�=FG3[ؿ��d*ZhSF��nf�?�s�K ��B��󃚭���q��#]��Y�����Mae����Mq�{��L�,�e�0 ��[�i%�7�i..��sO����ŭRl<�+���������\��Nh�K�:���@r@�k���C#@ҍ��--қ�( gr�8�$�9j�)x4�ky��.d�L>nQx�_}jY-Q@���#_OG.S�ǆ-ߜ[Ã��qin��ϐX����;6���[�$I&��as3���A{�����p�����/zK�^�~ի�{��؂l����bm��q�{�G��;��%Wu sWY�*r�yɬ�.4���^�8�[��rr-�I���M٤krE=��JjU��P�j�չ6|C�cZ�s��7����9��)�k�\���ʤ�3�w^���n�z)K�T5BR�]��N��?,��A�4E�0E�����L��q���8+@TZ8�a!��"� ��f�b�Ma���/����xe�MQ�6�$h����inF`��i�97A���24�8�I.Z%����(�9=wNy"�@�%�����D���#iI����_2���d��a��=�9�$�q*�L�u1�9���-�2�Gl�8���B��r��� ���o��!��AϞJ�ꧫ{/?\z	��Wxj��<(4�wJ�P�z�w+-Gh7Å�q�J��\�P	!]����Oa�m��S�@g�9&�Q�r�X�.&,��j^E�-Ѝ���Jj����潭)�@�S+�Sr#*Ќ�7�z��Jo�p^�y*�P�|�_M�Ũ\�k<jE����K-*hD�tܡ��0HL�{j��xQ��c0!VVq���%��Խ�_���$k�����K�����R�)�A�P}L�6l;|^�AA��7Vb���8r�8rM�[@�&Z��R^�Ȳ����$vH<�����Y�J~��Z��_��fo���l�߫Z�^�"Y��gMnII�	�OQ��뿕���r(�>��OD�u���
���֮D#���U]F3>t�'ܔ��ǩ���:��i��+6��պ`�I��Z�a#�췌9צ���(���O�������<6�4z�;�W��[7��Ә
����m��9���jG��E~#O�6�>��#�P��RaW9�o�SH�W��jBX�	 ��t�T���x��2.��`4Ϗr(=~�P	#�ݘ[u��
�0l)�\R���Cl	�dx�O�Ic4�T�b���NG�Zqi��s�����勮�5��+˱����ܨ7���������,gls)L�翮'���00Ҁ$�̓��]ѹ����ƌ�{&���^�����tq�b�g�5b�;��8���i��6w���@�����sd��!kjnzk�!h-.�;{��Y��;T`�����}���_�͒��Ď��7��h�,�� �e�^�&/������x��G�;Hb2�9$�3#z�����A��x0�zD��7����U�d'�_/�&��{��J�ĸ��.Q����L7���Ka��Z��沐z����P�N�ז�U&E
�֘�a�H�2 �-��vW���eY���G�������T�u����3L8���3O?���w�t����P�$�/��!��}((4O~�F�F�v��s8�3�G�o���8��]4�z���
,jL���oN×H �C<5�+-y+	R���/Q�/y)ǉ�u�l�g9M� ���?��n�G#׫�%��o����|D���5i�<�����*�geݚ� �!T�π�Q=tL�jߕ��Y(ҹQ�l?�<Soc4$3QC����*؟h�ʮ���-�P����TC�&���3M����{lp����SS~�E�	�2Q����-{�K]�%99�Hkr�s:���"^%W8�roz���,`Q�F�œ����X�:N�,tv|ܴ�$*R F[SK�
ӿ6�`x�[���rO����CC#9�4��#ؾ^�!/����`�w��=� ���$W<i�Hj8ݧ�t��<(/k��J��w��lJ)��,W��J�[�pf=+s�A/����&'e���N�� ��ۨm�B*�=��D٪�+�z�ȟ�">�i]1g�W������2�ysjsXd�S|���+��Gl
E��җ8�;r�c���ѐ὜��T�L�)V�}���iz�X7�(�%�PYa��[���v$M�x�vVw��by4$�n-���׵��Y{��������-��ԧ�����k_���ȡ�`�H���T��̸K�9Dc��x���/TD*I?0H�Z$�
υ
�:e��Rt���K���e�'B�r���b�w�����]�2�>��u�Jf&?�����J�
OFb����>���Nĸ� r�hgYk��J�9�heO7B��!�G ����".�������R>�
g��B����N���q�����#oz�*wظ�Y��f�r��7��}��O|�12 ��(�����	K�K����a.�bL�R��>۽���m}UsN�����E܌�ѣ��/9��1�找-�b�_��`J��O&>#�A;O�t1K~��|��}�1��͓#m�B������=�:�~�*n|�ᐧ�Z���4R���Ȥ�r`�-̟e�6��w��EL�5��us
?X���a�6i��Z� �7BsI33�|��*U���������SIdT;
��%�������^ˬ�}]����s��z�Pp��[4�N�������&�<p"�)Z7���lJ����ڎ7�v��u'�������E�T=I�Y��8����t'�V\�
Plj�H���L��SH*6Y�Vr��}���Ok�\Aa�?Q?i��b��V�H�}}C�}�H>ϢϬ���n�֩(�Ԧ��m���臰=HP�)3�����4l@�!(�X�O��|Kzp9(��j��_�}D�Z�AU�W�A_��F�S��p~p7(�w�jPnr��tz��i��Ԩ8kk0(��6�޳�VN���3�\��jm�GE�W�W�e��{cӭ#7$2P+*�P X}�$�$�YB1Ãw�\�`�.}��˳8q���ݗ./-�U�+z��A}�i�&Hn�׋�U�[��W�2}s�c
�d`�������;&������j��ۏ�RC.���Lgn�q��Z��9���%�X�����S��
��� �%��C�9#˵,ɕ�-ŀ��Cђ��HZIM�H�'�<��M�fC���������8�%ķ�),�~�#��`��+�F���虼8w�16���a��� l�:I
I�!̒z�e�j�;�z T�G���0f�F9��"ٽ���dd��?  c^j ЬW����dr�<���Ҽ������y=�+u k��ɿ�����"g�1�Օa��������`i�J@ j�ɚ�7�P	C
ɖ$fxXj!_q9u=�S��/ �uwZ(o����Atř�E�u�s���l]Kf���;�3&�m��<ww��78������[3�������`^C���s2N��Q�q�z۾��!���<��$O����7`��+�t����C(=���T:2�$x�/��S�j�[eC3O[�EN/�eGI� ��  +d��*���i-妝N��6���5�D�NE���q�[.x�XF�][:��
+�1���t���G�������;=F�pFj��g~.�i��z�;�3s�>�t�j�6��ru'�i��7��l���Ac��Q&C��Ҩo�ث�¾�&7���E$;�0���l����=�V���A�j����x�w���2�
�湪R�>!��t���&�1TG�[1G0�?	�s�6�`YF($��VA��x����H��1jԋ5ߛJIN�!��>Ѝ|�f��QTQ0[�8�f��[ "��%�*���F|5)�M��+�~�t�V��0�}�e��?Uoh�PC��>����f����B�DK���T��H�)%�!.��iE����=�j�&�������[�ᅰ�_�*��_ �~"����Rma�8����(㝀���,yq?�iC�@ĉ��j�����F�n�]��Q�N,��ȯ�ݕݱ�x��������Ϣr-��+�`��7��"��Ih��T{$��'�ޕd�!T�to�~��ҭu�'|���,��g�9��q����$���cx��L��j=K���/��Շ�±�rK��m�$H(}����1��)�K�_�s`��0�kp�>�8WJRI���_n����IAU��Ϣ�$�k�/(�)��i,�i���㌳�R���ѷ�^�8��J�Z�5�NvZ�2���=$jR�0�BT�n�<|��D� ���Mf+{�ǲ��|�ﾂ�RhA��
��	�Y=�2�#j0 �[%;�Ҥ���qK��6�zKO8�G���dJ��}q�����	�X㄂uGf̦�O�,�%� Ɍx�|<{1p�А-Z�������ݤ�A[d#h+�8�^��y�������o��R�C2��G|������FM��V�9~T2����T��&<�������vY���e�L���-��]�
&@F���1�j}�fK���ŗ[6���r1����K�����ͧL���%��8A���\�>�V	B#�nO&�W�F��������*�I��?��{ٗgJ́��lx���XَT��+m�զ�]���K�b�V����:���H�0ATd�[��Vv�zH�G��g���c)�jH��gD��B�dA�7uJ�j?T�
gW9���G�o0�����kRO��(���o�5�f��N�M��֭��I��~���w�x�����ⲋ�~��[�|<4���!�Ui=(��D���� �.��Uf<"����L̍��M���엜�Aޔ�%q�΃�I+���P��DA%�kY�I�3uvQ�Fz[%�
Ć�D��L���tw�p�\�u����9t��2{��V�ZBV_���lz�?�-�G��1�/w�.k��n��? �~R~��sߚV��V:s������ג�a��QZ
F�(���W
�5O=#F�Qo:�g
�0;�������:no�&o�Rů��ns-g�h�n�����Q��B)��)���w;�q�'��4e��c(�c�σN��0�Z|#&s�}^T[6k�L1���
Q]"p}�:�J#�g.�(w����1R��ʔ�!�h?vw8􀭣e|ce��0]�x�ta"|tF]�D����4�:�]s�2���UD&��[�1b!I@dK�a��,`	p�J���6��O6��&u~N�!� Χ�E��XW�&`������1�N�¼�8qmT'�:���j���� e��0�y�\�!�u��`�Sw�V�h�-ha:�u����C�}rv��N?�0^�C������>��&B�,�yKC��.���s��~
�Tm�N���Z�F��'�㛂x�.�+i*�1��ˬ{�-$~!�=��%¼N�<Θⲁ�e+��y�Q��'�������/ʸ��[9&O����8wWT��A%�Ӱf�T-���W6�n�B�踸{WW}����%�.i��u��+��tŔJ�	�H�n�-���:up<��|b����gT�Zku�m?'��餕�F���D��8E�)�����h���{�@^���E��됅�?��5lv�������)�q=�)o����ȝ	kɯ�4SeƦ(��b�P��$~2��: yibR�ֱ�14|���@O���|�b\b݇��}�|-L�Y��L[�A���X����1�U-�փ=6��� ���JX�>��w[�^��mzJ���1�-����^�"���gE�fB�'����Wc�<�1M��n����Hُ�%!v�D�tk-e��w"�1)^�<K�kPIᶟ�]�ӊ.DqSj��zx�=m֭�> GT�k�}wqf�����T����=�1��C������p��&����E$c�Z���q�qƚ�);p_ץ��6�I������T�t���p�!�Qw�gS�����=1 ��5�m�jg����*=��0�g�ڸ�'�1njc��(�c� U���z,Ȑ�@M�U=Jة!�<r��udlFE����qa0|.��
����g�w[�-b�zক�O��hK�N�/Uf�t���|NF���t��7���'Ya�"���Vu���\��IFU���:���8�er�����Q�bPd����ӊ5�#�[$�ht�"ک��|���'�GK1�����v�y�RJ�@��?~��Y6^�"�oQ�A��8�cU��[JP֠b�IIT��fE���L���t�I���%�M��;u鏼ZVёBJ#PdI���M�Z/B?Y7!���ˍᑱo����<��ʡ�Am�(��;�Q�y���sD[�����9���;Kg����ӷ .�!.�޳q����� ��3��e��a��e��%邍;�:mY˧e
��(���Isbh��o�͛�->�O�bUW�n@�������ڄ�>�~кg^��jP1��+�CF
����5%����rG�$� ���z���Q|���oL&�Ⱁ��x�S����T���0�b��H3Q��Q������}�g<���L:'��u��q��Yy�1=Z;/o/�쿈�
���+���
�ԁ�m��g���%*C���7j�$><
�:�k������D~=�:F d�D��ϳ���;��1�l�d����
��'��fW�J{��	�vH`�������mǀ+/:Ou�Y$q-�g|Z)Q�S�]q��gY��Ap��HvBk�M�tٚw�t�N6p��U�m�2P5�O�ۖ�x�xo���rG��##��n��&T���.��LP���*�w�h��c�%���ץSO^x;\��)��Y
G$���ݲ|�_�Y�������x!
%;^7x~ߟ�|��Oܕ�ټ�K��҂��^��I��n�d���t<HR�v%�'��H9�^��:�Lݭ�C0,����X7�q��|�w8F���Ci�D$�
��	��#��xU�������cz�0��_��~E�/x���V9&���q���
Q��_zB�z���{*bO��؈զ�]�E�cF���\iM���Q#jпEi�V[��2�r)�,�%��3\���ťT�L��lx�{���c� ���	�~���af��v���Ui�����Y�4�v]-ڀ~�����&�xo��=�JV�;�.�cO�FX�5�ׁ�7x���2�m\�J}�>3�_<]�;��_�x�O��屏�M�q��4��Ѩ�Ucz�hS����o�0y6�՚�����= ���y�DX�]����L@���zUmf��j��n��_[ʂ�z�27^t��ؔg�����Z-���v(��,5oyd^���!�'6_[�;�]*����d02zQ�/`2]�M!zn>pB�ןH�HW>YWa~�Kc�r8�i�͹;#͓k8�u����Α��C����<����J�*_6{�}���řiqo�ib�d��Hh����x�GwA2��^�s��;��<~�4U&
�[�����e�*Sg�yv���1+��!�=x���߄%��{ gi�_P�F�n}�V��Ĕ���e7g��k�������u������$hJ��/�t�}=�o(?(t��ڡg���E���K�a�N�Z�t{���*�1�j���0c[I�	Cy�`u4���x�,��YEO5�>b I2a�H��iO��;�����zqD�=̰b�2V��C^�����Z�s�%4w9S��}�O��7-m[d�4����L� \���F�lc��ǭP:\/�g�cAA2��=G�ZV_2w&1����!�o榻�[{5ed�b�&Q���?CN1�9�(�S8{ֈ�g;���.�`�ઑ�>1��F�����#��W[;�[%m_�q�EP�0P��7-����ñAү?��� `n(m�H�}�0#�������A�y��7�	�n�X	T�k�:/O�/�l���~��M�{oD;5�^%�qm,27����f^vP�j[���һt�f�ֆ�T�l�,��$|��v��k� !Q���'v�;m?��z+��R2��	d���',Q���%����6�%��FFv�x�_���-��%<s҃_��N�s�k��f�X̓��J��m�=Y�;~D̽+VI�`^3ل5�|�o�����[��;/��:�Q&AG�R9�T�_8���-kc_���G���G �ŋ��+��'$�,��x7��i�����!a�R�O2+%RA�2מGq�8���o�.F<"�5�<�7B�~!� k{�m6'�a���b@3�A�"����WE���Y��(R�ׯ���E��w�E�
)f4��t��U0���v穕�FEƧ�`��p\����Фi/�:`���#A5���*L�>jƉ��m������XN_�7$ |� )�-������t�M���^b@՜�z%$=D�ia	{�6B����X��W�̈́�����e�d��+X�jEm��VP���2\�(�a�{����暤j8���~N�A�>~�f����	y��̙���{8��k�/80u���WHC;���d(�q�V��g�nj���(�>�CD2�	��eP��S|o2�j
@u���çˉ"n�X���@���S�]��כ;j��z������.��7�8��k�jA������æO/o꟟?�Y9��a�zM�9X��݈��L8�GC�t�d��uJ��3�����������W&���ع�&b���f�ab��:�3&1����Äc��6����\���"^�h&��G@���6Vz���¯d<�|��y�޳���'���U>>�� ���9��F�a���pe������%g��ޅ�qb�U˧0�]��yS�.�]�}�]]�\��qy?
���V�%$2K�H S���o���!`8頎! �5��+���P���bO�������'�/��|Ѓbh��A�$K��p5���
�\��+h#��9ػ�VP��I[�qɆ�0r�O1�]/,�ܢ�l�T� 3���5]Η7ٳ`j/LpC<�B��`'�>�T�7��4��M	qC��Gm;�Mש[�d�4˴1�*o��L��MMv��Q���Jw�_ØEw���/��Q8��3���b��ga`���@7;���.��M({ߧ����`�����TP�U۷f�>aC�I>���"r�ʲ��\��B�,w]���Ϻ)."cU��O�%B�i��*�kj��8He�gG�"ny��ſ���v|N1��$s �Q�hX�x%Y�%�RE��!"�͍ bH0� �J'`��d�HO0B�����u��E��m�&35���WUT����/�sSsY��_\��u���.�F嗡�D�C@aEߋI�?3����dQ��4������5aU�ԏ��6�\�ҹ�e%6�fN�ǡ�}|6_	���R4���g1vq����OF`64Zr�3ʠ{V?~�hВ0Wey���C"�	�
ŀ5�A�_M�*k��x$�F��Yw��!{��A9����kg^���8�W͡JB�� 8{�nVn���H����%ˮ��"3+4��ٜI���HJ��o
$F�2��Z�		4fG��ae�s����U�\�������������%"��drY2e��;��<56n` �u�T�u�Wyj�v�Q>�g1x�9�V�6�X!X�:4�f���!QI��ŕ����|\ۉ7��E;��
r��ݢ����Ye�W~�ʩ)_^-+K`g�|��T���<#�#��.�1ѡ�Џ�YA�_B����j�M�u��V�t�8ۙ�]�;e��A��Q=�!|��@_G�����<gƴ_8]�����3?�`�d].e�����J���~�=:R?m2� y�m���A=UR>*`��Bn�Mi�A�M�d�p��uYkk�۰�}�����r����
�1Ln�N���׃~D2n���ȼ��隗=9e:61Lֵ�VZ(�!���r���Gb�꾷;�섔͍��5���W�f�U��+����sNv̶%�9!VޙqF�|�N��E�I���n����Zc�uq�����p�f�Q)��4,6���"ղn}�TLJF�/Yw>���k�S�d��3�Xs�&<-�&z�ɣi�hߎGI[�=���	��B�;t8�HN�f[�ԩ�	>']�Hv�G+���Q����`���(K~R�j���Ϲ��?�������^ux^�Y�<�  *�[g
�ux封 \��0T0�+d�R߁r�:��ϘF�oN׵s�ґi��瑕*��ȂZ��"�0Ӽ�2������ypVv�VΈ�z��<ſ�7��(c�gPM��O��3%/ҹ�|�����/Jl�m7�>��ǎ� �����2�*x��N�3�-��³0uG�D�3�F�l��[0\�Z �&c����ֽm���k���r�Ŵ��x)P��Z)��oS?&a'\�N8@�R����#�s�s2�é��Y���r�n�b4������)F�4H��h�Q�]g��>�h��j�dT|&`4�����yf��c���CN@
>F ��\+H�&�ۼ�Ƙ�ޫi""k6!��So�F�ȓy��e�\Դ�X\� #�E�O:[� #mD�����;�����̒��}�$��q�FgY~b���-`+�����؜�-�|ҥ����OWh��"Ya���!O-#�]c���E�L5.�N캵2�/�ݬ�T���?Z5��	�@��*92c��_!�� h;v�I��]��A���2n|��Z�Y�,�C'�}���þ9� <=�D�9�d�ͮ���J*�@v��A���6pvg��I��Z��d[&�=�ڵNj��_��s��
��3�Z�zp|L+n�^@M�Fl���ܦ՗�b�^���lV�U��?-Ǝ%�OC\?�+����g	M7 �h.�ن��/መ\�3�STL�u���`ґ�JT����S�H#����Z?���v����E�Q7��KڳٸYߝ�%����L7�݆ƑH!�!}\+�6��y]�I||�E�2]���f+�����T�w��}"��%���#J�k��n��������|�#�W:0f�irS��+|����>�(�Z��8�d���s2����bc(nB����8�.	�WǪ���j�2@FL��M\E�G�;0,C�d���,������T<���6��u_�j防;7{F�6]nF���j|F4��K&HvG9�9ڤ"*寊��͐ �ݕ_��Y6|x���o
v2��)�:�H1�s�X����vى-����jf�^�-��j~�Vs18>�� �S�C\��ia^Q��@�4g������|�-��F@�_7c�)"|^h�8*�"ll��*+uU�}{�Fm��\^"�1t�v��ț���[BX�qpY��)������6X*��>@�8K��#��o���:-�$Z�%TXĦ���r̂��C����Ǝ���//��H1��Y���̷rw
��9�|TDL7������;�����ڛ>��1����)4����K��[��s���f��LP�:��?W�|�$�~��k谦T������n��0Ƈ)ٛT���`^r+s镟5�/9J���m�++�7�^zs׍EE�"i�A!�k/F'
��;j��_m�$�\?s��,mdK�1L)��W�e^j#���zj[8B�w�)
�[I3� P��I�Iζ*iz�����\k@N"5�e����58���:��qVr��Sɥ�$��k����S�{������a��ރ�=����>}u� a�LӺ1�)*c���U*r���^��������һO�Ʋ�'��(8�rn���йD�V	s3��)��{�l�7�R�F~�v >y�[T�˿J٤.�f4<^7��
��Ƚ,��֟�K
e�;3v�T��/Z2�*F��!y^2����V)�E�G���mDٍ���hظQjx�'*�/�������e����}i}E�ŉ�9�ݟ(\R\2�o�.�Δr��d�quGZ�і[Y�|x�ڸJ���XPa�H-�<�Ʃ6����(P�y;f�nҰm+�%8���~�b��/�E#z�����$�����Z��}�(F�<�he�[��"�o�'��)r7{ee ۟ZO���T＇�$9'��M�,�g+���Q��el��Lx"��K;ro&�_%�@�U���"�(=x���:/b�G��U��j��h�,-�ӳ��#�!�V'���f+b�UϞ�0�����wq�Q-�7:���O�W|�_�z�?��]&1�:g)7��!z���{�$�9Ș�KW�m����7�M��,g��g.> �� yv�=B9qi'�<ɹ�i��ΖQ/=eQz�Ux�oZ$�߼ǹ��Z�H4�l��e�IN?h�e�j�w'����'ubB�LB	O��L��g	��f�����M����U��;������ţ��������<|����n����Wͅ¼�S��n�o\�a���m�鐒�8�ΫvG��O"Tډ���Crm�k`�uj�Um3��;�s�P��f��p0wH���4��x�"������Ӈ�R���a�xn���Tn��<��0S���yÑ��ezzKP���Z ���oC�˚e��rr��DDG݌a'*�>�ơ��7���O:A�"uk�e&�lg��Y��f-r�ѫSLi�{a4kĐ���K��P���* u��#��_�F�ȕ�;�-k�=�_��h	Z��d����l?U�m�bx2�Y�5\�T�5PƢ�N��q�� ���c�e��T�?֟@��������~;T^��D���j�����exw(�k��a�]����㿙&�E�*��1��KwfȊ��2?��7J��箉�6��,1#�en0R~��o�xe�o�O�c��"�3Gx����m�'����q�[��R��i�m�r�w�:���.ҩ��A��.���W۞�b�d
-�9�g',{���8�y0����@��ء�6'�����q�϶���a�%$��x))uQ�7�[��zp�6� ��P4�{V9�3k��5iudF�\x��n�|�g�[���:|��x"������1�N������
z��rMK<�F�f���W6��J��7ܪ�wK:�ծǼ�O*:E���pE;_Q��պH���p([�1���`�^�ZkuD�&���"s��~�!�},L���t4����<���K�%<��+ ���2/D�h�l��������u�0�@��$brJ8s�οڨ4��Y>`$C,r��O���!�R���,g��9�*>(��PP���ȷd���;?�����C��l�.̥�k���;_��Վn3�7�ڭLRb�5�V&˃?�C���@8`P|�J�v]�&���7��`�cy�!oxxms=H�*J�VH=��;Ϭd�ؤ�2k^ºT�@�~=tnͦ�����&��7�����q�tN29<�}��r+@�t�!#��9r~��m�y�>N���]�([�}W��SA�n�� ;����J�b�J���kZK\�J�g�G�[�[�Hp�T�u�?�f";W��4��T��[QGH�.�w=ަ�:d����`�HT�Gn.��dg�QZ�g�L1�Jve�^��m�[7���q�W�1�J��8�z�}L�
꛹�)���� "_"cir�CH�n۶
dP�	��d�t��QnfR�^v>��:�6��E^�*�`�'=��r;n+�g�Gr���Vŉa�ד2����L�^�ˣ�i.�'��l�����&��h�Xkp��)Q���fY���9������t�vI�)�oI6��W��6f�j�Ut�Lb/���E}���)$2;�15ݩ��~��qVN���L'�8���ۈ�3K%��"p3y��-�뗂��G�:�|�@.��l����=
��d�הV��n���+ |�D�%�R��u��Y�X ��B���<�7�¿�0�0������S�ky��ۦt�K�W�:\�����1�҉*�*}��v
z��1�L-�����B�l���P��сBB�L���(��ztŦŝ)�7��f��m~2�`���7������&NiԄ�Xq��gR�LۛC�.��&�:�p{�����Z�MJ��i���CiQ\��� K��_�?c$@�9�`r���vO=����9'�,�w���������D�~�!ӈ��I���?U�+�b.��4�����mN�����p��#�@>
;�tm@zB���|	
I��� �o�2�l�<r�5,hv�oHlk�M�z#������������Kb���
X%j������h���0y�j%��rTI`?��؋�aÂ�R"�Q͡�c1V�mJ�6-�g��@�[)<X-%����V�ufw����Z}Û���?�5~>ųRT�FWǗ��*b`�'G��wAn��q���0+�=�\a���_��j���?>��kg�xB�*tӭco]���[`� n���ۧ��w%1bC7�V�%����1G[�,�[�:�F�D��8{e�0�5��-���dC +<�*9�R��:ghC�/��
W����ʉ�Q"���J�j�8��|Y�-9]&��ʱ%�JkD��`�C$�V�ˑ������l8|��q���|t~z{��7�a�ARa��I �ۆ����H��(U��m�pX�0��?@�C��2I\��PV��rO� z	5*
&Ƴ�&ln�UR&6�a/P+�pߗZ$lH�hn�����r��s���D@2C��ij3�C�k�kh��ܑL���}m������y;��񟬻i_]5���̀�_�g�fn��.�C��q��X
�D䬝+�E=�\�36!3�~�,���I0j�����F0��{�+��0�����u6���{-�X�bL���LBP�#	��m���n{�,~�a9�j=�ě�%N8��?`���:����rR�� ���v�m�����8F��@�>Qi�v�-�q����u��ccA�^G�+��S+T���Zy�l��Z��*0O�%�����j�4��J�ŗ�U��_� ~!�F�r�(h�(3�z��{�U	@�%���ɷ��輷�_�ɋS��4�s�-�+�* >���Co哲�ː#m+&���Y����{/�ñ,��ݺp�Q�J���Y��+m���Y
G\ګ�]u�w���9C�Y��X��̚�We���䕚�6�������y���A�z��$��R��c)P���Sj��*�Se]�<�j�#�������ᛯ�y�,��>�EU�2q�ۤ��Nb�{ɿ��"�h<~D%8D�U��Tz
����c��_0�*��+:��g<�3x�Ae���+�?�N�j�M��J�͌/�.66�%� *�W���,�L��k&��u/��|=�EWc,��&������,W��dч�uE� �ă�� ����l�u�ZZh�EL��� v��a���4����\����7zS�ޯ��R�Ym#:'O>�׆�3�8hN{'m��Z�0���X똫��j� ������eel�j�c[a�Hŗ㍂ӄ�#��z:y�E���L�o�T:�7�&'!U��|�L��|��a�op<"�4T�j:9I�y���M\��S:�Ӯ�3Ǽ
1���܃������1C�w}�&G-|�iL�]f�?R}�O��:���tOx�&\5�ү���ǋ�ѷ��]�D��4�qs��6�KW�c!�����	Ј����F�)�ZG�����Jo��Zh�ɱ��B�r����HRD �0�i��C�A�#<�B�w�A�ߵO�8e�q���	��ڕ���O�"�s��Ug�\F�y����Qn�O'����46��f2�CRk�C��*�VA����C>��,���RAR�ֿ�;���Gr�(#��I�Ҧ��&E����W팮V+[Z����>০��b���I{�M�U��p�e*Q��A��wiK�1k�-"X@j�M�ԻZ�Z+H��3l1}��6��=RTf�}Ã#_����b�`�X���X)�A�E�:�rl��r8�빙�J����]6����q}�"z-��ۙ�~������j��hO0-�O��2DU�����n(�2��%�T�r��k?����(�#��ÚU�h��oT��D?�8���n�m��k�0�i��	"�g��5���N���ҙ@&'p�� b^(������gɉ��[�G�'\�CIkp'd)U����?%��[SX�)O>�C�j3��Lv���A�G	6I��߿kp��N�)
'k��7����&�C��19Z�y���1_&W>iXK�r�A��$������e��kjc�����G�%rM\����9�;	)�4���"Z!U#�%���m��M!�]E�Ḭ���.x���&���������=�:��j-�`eޝE� �Ǿ����E'���
��'���$�Q`��ެl�N��9x�������t�������m�f��s��%�0��D�f=�]�7��(L�a��{)�jWv��O $l{�s��A��|:�8A�M���g�^��j��`;���yk捱~�4�[�>�mxQj�f��Ԅ��-#!�2$hq�+�j���"����^�r^����<�Lɖ�
�����:>�AKC)WH���E�+�������(S���xg��7V�=��#=�99�hС��U͟�+������=1[��3h�ߺ}�_�z���B~�==?�z� �oU0�v��<�f���+a��̫��r�0u�98��_魍v��Q`л7���
-,�f|uL�gϓ�(k��U!jXⰽ���s�Vl�OZ����0h�����<+%h�����yx#��,a��
Ȧ潸��H�6��p�r�E�U��y1�a=����Vo�5����Ĩt�q�k⯕�c�R�}�,��i�5����cQ<��0}�2g��+*f!�  A -��6���3����t�ѻ~����آOͤzI���"5��_:��0�U5�t����E8�x�|q���6�g��dUQ��b5�����U��f}��?}���"�j\�Y0q�h��põ�Rc��t�pa�#�*e��	����]6�k��-������3��L�Hn�3dS��Ѝ��]�*�pM���6K��"Tq7dC�P�o�%>��ľwY�և?VT��� �\r��+C���`РA�d�T��0�5y���#b�0��(�u ^:RIY4��x�),�ƕ�iUG�rJ����2��qznH���@�ܵ���K�%ّ\kýpR�4ۊcC����;azqW���Ϸ�*B��glE��a�ܾ��"����s���7��{�[��g�E��hR��y�ݶ}�G�9���=�>R��Fo�L����5~ �$9����L���[�vr��j�Ĵԓ�f�Lm�����,p��������f�	'Ѡˏ�PNZ �>|$�)�8m��*q_v�m?l_��N���p�;��z�o�^3S��jy���{�\�K�N�l�'w'�~%����Ω�/�@�$�]�E��nb`+�����ݢjy�4�k�|�4�C<�� ��I� d��o�ă����6n�eT��(��*?ن^LF�T�w�)9*���X��E���$Ȍ-���K��(];��5>�ҮzT`myIp
�[]���"_�r*���ĭ�m���þ"�ʯb`]�a�>�ضU_�4*R�N>��tQ������aԃ%q����2��УA�u��g�y�{�M��)]�O�Z�Ͻ&�I��,�3E�]<]-�l�b[
K���+j�x�9� ���1�e�e��0�V��c��:P�[Z���=�����}���nR*KL�F�MS�5������=
�S	e��>��-�n@+���c����_���ԅ�ZR#������;�j9/�<���Ċ!�s��֔�
wn��F2��ͷS�z��n^4<W��$���1�.��`�ו�a�r��	�7՛Y�j��ó�G��-xMڏ��l�rpW��["A�z1�� M��L�zy7(!X��β�	��+�JM[�u(��;����#UۃN��-��F��i�l6E-�z[!]��t1��1DH�O�eE�L,|���`��id|�iV錦QW���i<줜#>+� ���;t�{c!��xc�	��w3u	�Om�"A�H����U��]v��c�ا�-��W�L�>�&�SD���<4���1ǸR�M�9P0�����1}U���E��[�Z�Ҷ�,-��Q�C� DM��j��vؐn�Y���j��Y���%[�h������
Zs�CȼK@#�졗���=,a
F͑*�b�>��$0j�����E�b2�;�㛀�F& �Z�r:��|Ο�K��Y����g`.��^2O�f���o@`x!D�1��λS������D}n�V.�3�oap'��^u�=yBuժX�l�>$I	�_�{�����D"͟�U�����
�j�"���;���]�aT��T*���d_����B݃�}��tq2u	�J�^�:D5�A�3�!�$c[�±�lO��h�Rn�h��v?��s��S�E�%5�p���8~"S@S�l�d4�^�.|�����q��,?��"C3CĂebY���"�R�,�m�q�ݩ-ԝ��K/2�~�R���1{��i8�l7�r�)n�k��"+���v,Ip8�@���W��.�I�ٮ ׸�wF� z�	�Oʪ��9R"�� �mك\�'
_ڶK=���j�͊���>�'��+r��~\pk8���?'�b5C���DL�6Y��b��4�B�p,p����m�A<Ύ��ԉ�[�@���~F yp�բ C4��X�~���;a�Z���Z��#߽� .�#��m�xN���Ȥ�^(�����N'ژb Ęڶ��ǅ��95$���N!{Ԇ� ����\Q��L�-���^LQ�K����r��_K�Zk���L=���ĩ�*��������0%��b#Q���q�Y>$��""Wz�&�>��4�n�xy�ӋT�k��L���>Jǿ�F�Q�?�;TYס~WՔ�zsb���J,g|3��b�E\\�\�C�'���՛�r��xb��O�)	�Hы���X��ѐLr����T?}�+"��.���_cz_I���el��p_+��vi�*�(��G�Ér��8�4��q2F���e�.�F�h�a���x_��L��" �v�(����:�s0�BÖ��7����o��3�.������J@��oiA��iJ������%s�
*�>$c?��8#�'�h[��a�g��(��rV�J��=(_�T���RUR�)XA�;3�z�����͟v�F�&�#����:�o�k|.��q���4߬sT����
@��c3�@��5W�fA��/��mǍ3����А
���#�ű�H��w���u��%�m�"I���e�3=uޠZ���g�{�~��xD��E�WǏ�V[h�G�eY�d
3v�t���-�� E� I�}w8��ߘ�����z��&�K]c�+ʨ|.KȲ�0쐭�����i��������^	;n�M��2R���gRѴ�� ���@_k�*A	Z�_���/�E��@���e��8K�W6|�P�w�
(�����z��9�-�䪺�s���>�e�Rv/�e������o:+�
�."����mA]�jO(e�̐��;7���,R�����d$ܙ��v�1��o�xZ�kFt�@�`+(��cc�bHl�!! ʊ,�E�7���?�h2b��0=úhV���ŏ�7�Koa�&�R��g�q���ē�/=ʉzJ�u5P�V���ܘl�0�o��5�c��V�8?x{�i)��
+�H�B���9�>Fy)�K݆Zs��}�$9	R@�&��_�.61�Ҫk�Z�ai��#q��z'R�Hc�ɞu}�zxX�B|�	+R�U���Ԃ!Ҷ=�k~��Wȳ��ƹQEp��?U�˛���L�g�w7T�R�eM��ekp��.1�8�K���Y�ŀ;���c�<�2[�I�>s����s�����Z�o�
���ƒ�Ա�V��!<�8�S����`�v�����q� �[2#;4�Z��m����D;��}C!&�7Pk;R�jh�=���!a<՝	�¡�2�������9�4#����&��L+�����|��V�bO�X�Z*�3���f8G�K�w�k=G.;����l�`H(d�ߗdM�#+��uA��h
�n�d�{��6�`��L�m�&�b������%���.�D
��m��Z��o`��o�7{�3��'r�ǻη�F�7��%��sso�L�ڞ��3����E�E\�7��+	���z�
� �:��{�{�u��]��~Բ}��,�I��F��,rՃ���pq���Wo�W9~.~��p��h�,7b�g���U�m�}��hQ��l����g�X&����whb�����ǭ0������;�+����"�;�/g#h���I�;��:�3�YK�I�}�Q�jj��h�e����=P���!!���iK��]�o�3�?�P�^�+�UK��8���.��9��ն�����pź�%b��%���5G��(4%g����ʌ�#����9�� ¸��yM-�8��2��z���Xm��r�-��<����X)�Eg��Zz�,u޼B�tT���̳T5<|)�$���0���@́�nk!���b�G�_�dq��^6�
��;O��g�U2(���	�7(ū�0�KJѬ�9j���S�ciԒkl���\;��o�
��+��xׯaZz�s*a���EZW\�d(Q�;T��	�E��I¦!{�I�������V2�ӚQ�����]���X#;��QN�Hy��ڱ�#a{d�~ٟޭ@!�h\z]D@
T���8�-e_3��sr|�P�\�-�+��*�/AN1��|va�r���ڒ��4Qp+�����Ֆs;;;���t󌫤�7�*����j�g_������|������$����T�
nAy��\[��C`9�N�!캨0�qM�2��u��nI�ÊM<��.{a�d��ʛJ�cDd%!��n��,�ʱv]���['�{%7P�H���bC_�k�WBfY�k��(vѽ�{���)ɩd�_L��RrT��n�	5^�م»o�vUA��cה�Oۏ�z$�e�J�y.Ss���w��P�����bl�fI&�Jdfy0����Qr�@h��ג�Z�,1�"6`��q�ȓ�,�#1%�ц��
:��uL��O6�e��*r�C���9���{��x؏�5����Z�)�����H4*��yJi�D�e��^
f����[�P�<����-��cj���"At�}���6
!J���*���(#����"�	{��p�����p���|�>WpώXn~���b�&��l�z��6ޚ3�(O8�Y=��N��h�y&�*r�S�@��O�#��@A�M�&���@W�LX��DL���F,S"/���������˺�N����r��7��4gzR5�&�5�V۩�M��������K��-z�G�y.������P�{���$�\f���5	{o�)I_�aE�I�o�����i�[�j_\�����9��N�:X�A�*�3L}x��݁%��UY�wS�Ew���u�>��p_�?��9�n>yP�|`���gMXO/���kaؠ��c�ٕ	�?�|�R�{-h�����NT*Z$�or�3oԨ�el}\��r�S�'�t9!_�4��M�E\ՙW�F�}�Ѥ��� ��~.\��zA!=+�O}�^�Z�ǁ�m{��}���iJ�'R�hv������K�����E���eG^~K�����.����J��B�呅\�)�5%���UۉIj�.��$=�=2�м�s!�����R�V
��]&D��:i�������U K0bڱ_oD%����J��
����<�6��5��cz"3cVB#� �/ŋu&*���me�p6ٟf%�l�n�(�ߡm���#������ӟ�A�'ߌA�6�����\��u�G8gv^�xR��M�ٸvwW��]m�m�s�XbK�w���u�K�lV�^h��7A�:"�)B�0�d��~''��@�F�&�w_f�7\�6�'�"�	�hZ�p��%?�Q=6�R�.�{EA,����;p߅-����[i���J^��(����������d��2�!��t�HT��cR���4�#"��� ��u��>�v��]YhXR86/�[��D&/A�3�"�%6����pR�ǜ��]�?�Qw��w�b�T�gucZ_�Ɂ�4�Y2�w��4^���DL�*q� <kT������!v93����YX�n�/Xqf�닲��?�a�ueC3�1�����ݕ\����,���Ø����XIF�ָ��bA�9?�c���|�=r�W3qa�FA�E������w��l�����{�F���g�pM\f��jY��R��Rv��6��X�n���u��e7?�*�"q�ҙ�����ys8�I*e{�侻�GhF�=��QO�X�vẸ�Jٵ���3���v/Y���s�U$h]��#�r$b�n��B�3$)�@�E���Y'_A����i'j �)����ߒ�E�mB�y�|��q.��
�0o�,A��������y��Л ��_��)�J,,��}�����͌�0�?��Cej��([[2W�=�g�� Pw��r20��1����;n�q��T�*^k�X�u"(J}Ƙ�_�/ɘ����o����y��sg!�V�ڿ��c��ȕ���<a�Y}���{!괍wܫP��b)pC�ï���hҎ��9.:n��3�$����$�֓��Q��Z�X	�c��[����d�>�n�{�b	Gw��8�B�r�(�3h<3<1�N��r�a�ym_���HJ%#qf~'B�=G��xg�^R��;#@}���;m7AO�~�s]��~�W�W�e�^2���'C���oXp�N��N�	RAlyA���������p�*R!Ov<�.�r�#�ұ!��هwQ�J�R�K����B������t7<��(�&�ھ.�0o]��m�:�)�
� ��a�%d��!s�4O�6�?B�3W(��$nB��'����ѩ"�0�;�ڷ`7��o5����A�j<{�^�1�F_.%��v�?|O)�d�
��?Lqn�J,4�z��9o�xyԊt^�Ջ��#���#7l��5���d�f���.��j�K����w�Op�h�2�i*ۆj nb��M�!�9(�>d������+t%��smu5vc�qA5U/D<������H�c�i�H8<��� ~#�3��w�V��[����6�!˶�pT�Y.��`-�P���W�M��|ߢgleJ����0��
���A��i�-˷Km�O�0�{�i��_o���l7kH��#,��mZW��ݠp���xz%g���{�i��Ȗ|���{�5�Py���#���'��G�DC"�Ǹ=;�<@[�L�ɉC;�F^q�6�A����|�闺wp��>-��ÓRkU3�vr��DF���I�$��,�2��؜���VO��B�b�fFg
�}��>e����ƢZ�C�A���C��aN�Af$C}d
�7fL�߀�V�c�]1k���"��}p��M�D^�(�_E(tֱ�'j9fyo!Def^�,��[�.��;�ɂҘ���OUƏ�b������j��*��Z�b������U��ԏ'��6o+�M *<��L�G�;�6~�Ts�m�[)����@\�i�$Rܲ�!��
�ݴ��O1<v\����;�wO8�[��;Vw�Ԣx��I�wό[�x���[��L_��wÍ�#�r�C�G7H� ����f����x��Rr�$�
�;���&;}z'-�������Ir�LuqAe8��[4�HQߎ?��#=��G0�%������X�K��
+���ɇ�2�;�5I���u��VL��1�w�2�e�Y��/��=��?=MNL J��Ge�L!��bY�
:f��D�����@�ُ'������,���Yh�A�g����~_B��ح]���3����J]�\�.�z��<,��Z������e���́������e�2�u�Q�U�^�Qu�A�\�{gR2S��+���L�: 
�I.�4�����>�~�D�N5��i�!o�;~�h��-?����_�[�Z�.��v�c⢬�۫�N_�t5O�~o.�:��g8N���+���yD���	v�9�,�Br��"��H��zy_�/�b��ٴy�y��r.�۵(qY�T�]p��_f�J`�s�Da~6�am����H��*�I��G�8M�UJ6&HM=7o�M��X��~8�`�)�a>����(�TNJ��DXYt��~^��֍�o�D��o�����}RTU�6�x$�Ǡu���&�������{H"K�۞ ��@�3��'�u=J�Rvm2꘶-�/��}|����G+��suI���l�3��Tp��$JZi���Ȱ���&�#3�/}����o��r���:�-�fe�m6bǿM�	���[B��ǈ�	����aa��>�4BC��K�YF��(�
d��k{
���o _}��\����w۪�������ރxa߳��V ������A�	� �n��fZj愺�V�S�h�P�����y06/�'��L��v3��fo�h"A;C��V��\��� 3a䪾������q�sO�C����i��	��6
�[�B�:
Eh��w����Q-�g�Tn�#~���u0��i��;f^_���Ǚ��|�����x�-���,&1 v��@ܳ�%�P05Ջ&XgvP��Y��8�
F��i&_#3=܁�P���*>��|4�-�)-�J�F�R"�&{�
>�]�PD�T:�qX�����0��+��PV����1�[�3�%��u�g6C����y�.�
͑�U@����GZ��:�a	��q��?�f�&r~Y�'�EP��e�Um?.�bv�Gt�-��L\�o'�n�[�9C��.��!?�3zos�e�M��/���M��=�콦�
�)0n邾B�q3C3�ۚf���.���E�>��W���z3�j��d�m�gk?�|�K�#�f����m�&�?�r3��v�ƤW%���l_*i��'��˵�RJ�&=�r� �t�]u+����R=���8u|�81Fo��'V3ɺ��s�U)Q��R��>˗R��������^4͸S�}��<����a�ˋLX�.�m������JwF\�l�H:(�=��ijP.f7�_��ᾑ\Z$�Cۃ�m�h��;��EB|�2�=Bs��8X�MBtT"�kR�l�d�خ���p1��PѴU��
2l��\��|������4G�e�����⦀�>�!�P�V^��}���]��aF3y_����V6��0��O��@���[��h���� y2��H?�B����_������|��WPg����`��f��5�H��fG�+��d*�74��-B���53�ɡ:Y}�7���x��A����e6.��1?i�ݥ����)-q���
�a�D��EoA����h�Ϟ���R:�<��MoZ��'L��;���񵦂у�9����o�/�]`�����Pel]Q�$>�T�8���L^����o�-Ua�$�!�ҫ��ؽ%n��ҧJ���p�{��ɪ8mEB,�!U�T�-gm�xb�l��wË�R���B��O|�Wz�/L�!;;_zn~�1>�����c���K* �����u�����Ú��H�]x>�B��!˅e껈����Q�/�"&񹖍ny�d~�`SX"��e��7>�/�Ҡ=��~��|����@�H�d͜��򴖤��xs�q$�[{���&ҵiBY����ԅ��»�&�ͦ�2�K|扁b7+�:,$��<
�>X�Qlퟋ(�_C=�h�h�̾�g\���t�@Zڢ�^!BP�A��w� ��\���"z;1o��tD������)������=�3z�TV��,�x�eD;�������%7��qjs�J�D���\���YjG/�0�c�CZk�n�����|0���K�Q���������`��;�}�	���E��nƘ�_?t�Ad	���8l��q��<��xC-8�ᳮi0���(��e���B��҂�Ҷq'��얐&�1�F�3��]��9���f��O��;K
��"l>ri���@'��x:Fi�������ζ���*%{%2VoM�Ǿ�I����R�p����wZ��yY]ϣԤ-��=�	�� *z��/yɶ��� i2@ؼ���P6��ۙu��/�;\[��x���|V��|�Bf���9�J���E�&���*��*��V���q:�i���:REzD�i%�����{2�W�AN�[���Cݜ��i�E��h�2���N	�G�6ux(�tk�;�,N��|>����~Ý�F�bE�줕˧�\�Kr�-��mc.���S�eK�����p�����7*�@��#[�~&�h�Ӏ6����gu"��UV��O�rtը��_���
�#��{}�  �9���gJ���Ye���MnH	�(6�	���y��Oj�\�31�u�M��#�MP�W��tj`3��G\~�U����y����p�f�e�D1�T	�(�P�E� i��\>�6mZɪ�9�z��-=�`,��N���]�`t@=��	�b9��JvH���q���{��<�'|$��&ϐ��N{����5G�E����2�w�i�X��3"	F���t�3�n���{�"A�_G#g�̇�@!(w������Q�U��< [^x@��q�nm{���*�{�;c=��ae-R�:L��(�ݲ�˼瑐�D��o��S���2p�D�%�P�	T�Ҧ��]O��!/A�C<$P�@��o��0���TL� <(.w誙��FB��>��+2����@R�9Jt楂8eJ9����܄�kv0&�ոkJCdy�p�܊B%^g�Pɭ1�/����l$I��<��[i�\@�7v����Uß�~))s����%Mf��f�&�@����i��� �9���z�/����[�	20�d��CӃ�3aM�W�ě�hc�V�����TY�\�pZu��ʏpc�oހ+�a4feg�ŋCv l� q$:sa�1vPU�[C��2	�w�ߊ���b�lPZ�?��ݼ�2�N��4�.��L�v#���H�������-���6d�̘���j5���JP�+tv!��mOu����.s���Q�-Ewm�U��N�g����(��Y?��z���?!*���ly�4Tu�?y��LҦ��;IU�b__�:� ���0��t���ܲ���	@���~�b<��T�\� o�o��2�4�w�\�C�7��љD$�$���$��˿�콴�PD�	��::�S������Vc]?�*�ϒ���H ��(�=�b HÞ��-��7�5"Q�QQ�
p�|Ap�����<zH·�1�YG�MAD�z�@Εr�;�e���ƫ�&��_��r��Hq���<\��&�*���_h��~��<O�/DW�n�9��s�Tfv��/]��0
=��5�����#������R�Ԡ�_w@��O���u�q����q�s���Ǻ�uܸNT{ܩ�M��rX�:PEp�
R��v��T�3��Dqc�Eh��]���-�R����;[4j#~A3ֹ|��5ѪNTw2�az�﾿�v�y�)������`��-���;��~^�F��RFd1��MO�g�o��^&���,R ���$�tK �w�& ��5m���gt .��Ҷo"|�Q�h\�4�Z�~B��a��k�r(L̀� �u���E��%�=� �p�Ї�N��H^�<��m�z A�퉗�v4r^��}��Db�5 � �5T�_~FG,-�_7i2��@O�|G"�0z��S�Q~9(�v�4M���=Om6��3j���;� $|j")��w��5K˪r���E_�Q;�;(�V�����zk�t����Rm��.�񤫱Մ�5�I�9��`�6�Z~�N�mqY����:�Y�U�N�;� �X�k��!WI�Ȑ�e�>o1ӟu�����]d�=�6�~S9j��n�"ᳮ�r�� ��f���QM��ɍ�ì�3X�N�_O��ۇ�Q�mP�G�$��2��\�lL&�km��i� 
���YZZ��JD�
-�(��R�T������7V�Pi��/�\	��%cr7v��nL��&�c�~��6@H�S�K�H# �`s!�Cv���XE'�/h-P������� 3&�:�F�+̑����Ճ&t�-}>��q7ͭ�}ּ�V�;n�X�:�W.�