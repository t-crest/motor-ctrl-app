��/  �~I�⑵�ۥ���"�\�ӪI���%��t��]l�:;�|P�7�|-:p�#�tS�����H�Y��j}':�1ކ/�F:�d�ǈQaz͆���b9k��wd�if����p]s������W�c���n{0n��#��J�����U�K �l��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<��G�y�F��j��G�9���co3������m��_ȥ��7��G��h@���\��̩-g��l,B������w��R!�����Iy�5n|L��� ?�R����B$Y	v�b1=��2�d����������RL	T�$��?cM>!R	��^b��y+w���M|�K�\u��������En���^�֍X.�ũ���G� ix�[��ʒIg�<#g8%@y5����jܦ�8�a�=	��&[�t���h})B�0.�9D��Q��a��3V+�⤌Z�9lHAF/��c|7�pH��ARq�o7�A��K	Ѯ�w/a�����7Q��uh��榛��RS�m2f�##N��9>xLN��B/+[B�{6n{V�	����|���ுSCR��L_Bb�7˫@&~5D��z�_q��j�	�^�l��B7|�A����!�(GT �B�} �an�N���O��+�R�I�@�1��\�ߺ�qs�|!�:�f��5�4���Ŕ�;f>��_�ϪbB٧�ze
J����1V��D7��Ȏ�>=�<�3�����}���I@Z�>�o��t������s�co�� ���)�x�*������t�U�+�y�R�Xz8J���Vn�=_�]<�� ��»0wu#��HJ0֨K���z_ʆ+�J�Z�>G�J�
��*%a����!�.�.�?i=4�h(�_y��]���B��4�(�Ș;�Ng� 'Τ�f<��x�iJY�m\4�B� #~��-M��hoyt�Y��n��G�Q��wW$����X��H�;��v ��Ay�%�����5��%�Õ�-����~J�L
�r��6ɽc���|]Y=I�ӘN���V4����l7>��Uy�s!���hnWA���#��i?�:j���ѝzv sƞ2�l.˺吵��4�s���!� �8�^�(��M�x��e`�wP��}��>/�-Ҋ��w�M$U��@��t�c�_��}R>$�>�"�W�D{��kJ��`�;��RW�rQ� �i�Gsҍ|��~E��&���Ҥ���3(o41��"P�9����+�r�Z��yF2��/���H�*�-�#f�?>d(79�Sl���y���s�&ң�[���ԿR�P�T!��2��c �Q��c"��Xx{-�9DB���r�"����g3~1C�m
���E1Ն͑�!l�)���oW�?������D����l��T�-���<�h�t�`����V��p�\�G�E���Q"�ϭ#�����s+� G3O94�Z�V;P���c�/K�,�d�o�$$�8w#%�4�n���I,nr�>W�2��	�.�ɨ8ف:
���G?��M�V�=���B��4dS<,�TP�y��\ք�>l�C�S��\���uYڏ��<��^@��BF��;L4*�ǆn$
�%��J1� ӹ�ü)i���;�m�uh�
n�t*���O�nݗe���aE>����DY���]�|�}�DL7�T�1Ӏ�Y~$Sh���z����=%B��r�R1+��R�n��a���-^SJ�)0wWW�9;Ra� n�f���B���q�4�r�P`���~FV�X%�7䢺�6i�j����S)�?�L	�l.���6�ժ.S͈�Ni])���!�o�����J!� ������cs�,
��;��w8���Fp�:���cP1a+����'I�z� 4u�����`�ּOl�'�g|�;�B��e�Ŗ�ҪI��V69�y�af�b����<O,�˂��B2)����H٥�2?x�Y�l�V�;���}��J�מw�a�R��Y�h.�muەVc16�)\I�c����H�XW��+�����\ͨ���P#�# �tW�y��B�3�)�0������YG*^`�*���p�ٮ_���t�t�.�d�Ȋ<�*u�%G��zյ�;�S�4鮖ϢF��{����x�f��@�]��שDWf����	xl�m�u@��z���n����Td1��Ï�2�+�"��5$@~����z]�R��V*w7n�껭���	
��.���������bn�))f@
G0��L3�9�:�i}�E�9����:���|ط����1�܆C�dԛ.�8�YVD�u������[�T�PJz3I��	z��3��׏M��4Q�c�C9�4~��OB.��Fpy։����"��G\JJ8܇���7��wG{:mV|ܴ�W\c�_ ���j���8z ���'ϼ)� ���a�5=�d��N noEP�R#a�!UgФ�_��Z��`~�O�484O�:������ U����a�?v�&�
���K���,�'����}���!	]Q`��nM�tCҤ�o�ގ�&}���,z��|�D�-�,��M�t�(���M`�-�����+p�J��ѻ�].����	J�}��-r�)O"�����,'I9��	J��<��/��C%C��F!_`���)e.~��û�u����0�vڎ��󗖭��?$0��xm��]\�U7K߂��c�m
	W�μ}�d1H�����E���h+/�"x�`��߮������l�%g�}��_ 4�_����_'�c+��r�����n��K���U�~�aV�啡	|=Z�	S8��Η��:Wg�������-�ؗ�	@=#��e�jC������Q2���)�狐}X4S~���lu���T��͛������E������}��_�M���)B��Ҍ���}�%<�[q�"�ڃ.N$"A/����P9{�5&=��-(Lh�T��&���Ϫ�i6�N?g�a���@i�3�����%�L����|��N&��F��F���(��#u��Nm���G��
���T��m8��<o���Зl���#�ڰ���x�X��k�����LXb��3BơP�&쪗���'bx�=8U��9�#rAV{�S��.�]6��#A�}��W���~ ��G��

�I��lr�����f�0����b~#���AtT���?(�r��劻��
+<׈x�$�x�p΁�ј�߼V8�pol�?��Q�L�=5b :̌����8 .��(�gn�KD��w��#��.�1��u ��Ua��Yl�'le�dJL�.����1�V�X1�7���0���}ʥɩ��΋��K B~�Lw�g�؄_���7��2Bl���Dx%e�"m� ԍ�S��-eN�7Օ�ɳ:��rkUv&����-��o<ۤ1�2�U��F�*;������&��`��l�Tw���j.xho�$�Id>Xꑷx޼��Q6K<���`��=�M��� �#b���Y:_�&ﭒ]1Ny���