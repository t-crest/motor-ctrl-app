��/  ��\H�,��^h�1��&v��e�v5�GyVcaÙ�9a.�_�L�p�|����7�]{�{h�3�B�F�`���Qi�#�uM~Aacp�"��:�j�����zMY���)�&����%�t�9���^�ސ��"0�Ц"`C�j���P�� l/u�(��]j�^��<�J	9�yI۴�:Sހ?�!��mbH3.��^;�b1�A��Y�Ǹڢ�n��0-��$I-|��:t�	l�-��>}�2��C��$"QFyC�qp{d�Ǒ,Y)���Fg���2���g��}�2-���H�S��Ԁ8��x�{�J�c����QP��}���m�Q�xx,(f;�G��wQ�\�zu9鄁ntpi��z�|r���[l����)�/��<��-�έ�'�8�g*�fs�H҆��'s[8�G���:>㲨�ֈ���#lJQ������WZ(�b+�KJ�8N((R
�����x�5A	��3>�7�Q���`9��Iɑ�����ѯv�/���Y� ��঑[�[t�EH�ݺX�s�*��G���;g�Qʘ����/o�<�Ǻz�����n��]w���ӛ7�ɛ�@t`�H=Ъ���l�y{L�)�(y�.��l8ٞ(Ö����D�k��!�-��n������A;��ʾ� ��Z�֛��ݼ@ȭ�>W�:*���x?�xk�R�#ܴ����Lx��R2Lp���l�W݋���j
3�3Y��,�NMhF�$y$kk�M5�wt��0ӳ�w����i_��J�Ҍ�u��x4�'!b�ګSb����! |��L\a�8K�ؖZ�}��L~�;�L�������j��D������8�*��ȴ+�+D���nq���'M��f�
�"
��V�qW�H�X���?�qx�$eڲc��g���m�`�e����ēm���`��nĳ���?�870���}�윤8��S�������]M�k��^%#A �գɛ|��SD]Ԩu�6�n&���U��_ŗ��S&"�dT���u�u7J����R:<�w���w��B����L��|Z5bPct'�f�����GW����9�����]�u�6D+���Jl��JƔ� ��AJeS��C�r/�����.�`Uaq.tc�lBE���*�RyC�Z�}��gw����r[���C�	ߙ�@w�~�	\{�Ww�2��:̫r.��XF
hʼ���A����?��s�O���$x��`c0Kp7o_�h��I��u�O���uvүX9��!Ce��� ����� 	$-�(&���d��)��\���w�d[t��y�<1K���2��M���gQt3-�-�/��UW�+��e0�i8�����E=�W�B�M�[ ���x��*'�ĕ�dɿ�"�%khh8U:�)F�����"Um2�n