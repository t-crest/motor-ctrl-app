��/  ���K�;,�vS+B~r6�h���y��`ὩkO'�&ց� �<]%��7%��Y:���S�?�H�o<Eb�	����$�xf��S4���t6P���2���䫪^����H��:��.����gS����,D'������E��Ym]X��x��	��9jR>��6-롐K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!����ıL	���dG׉:�v�&7^ș��+�W1���_� ��Paj�u5�����Q��ߝN!(�F�C�R�������O$�����W9��	-�KT8q'�J��ل�)�\��Κ	U����VM��'(n=y
�ܡ�T�h�"@=֔�/q����=w�K5�@�ǻ�U�̅�/���1�I��P���D��!��]�1c��V�����4 Y��6�rrF�Ex���F�TT���&6l�'�c��~�ɞ�	��S��E���v��
s|gU�dG��7����d=y�]�D�h�/���a�2*���l��r$���9�vta��@3�!�Q��Nl����4J����{^"�{0IQb���̽���T�S̡c�r�5sޞ��x����B���d��S௒"�Ko͞����U������@�<|��a��
���PV�y��B
׸J0G� v��ʗ1�������H������'����<��)���H^��G�Nll�L����b�Β1�d*|��s��":'�I�R����?�M[��߮mě�Ƅ8=�H�>�r�.@=*�ɨd���)��5<̛�؆&��B¿$(�_.�����,z��}!����CU9�rL�A��N� ϝ��kt�9��, �	�9���%X�DK��Xt9ON�\�?��t��&�*e5R҅�����@�H�$��]Wg��w1���|� �ۓ%�#���PW:,��w��@9�,�ҷ�������,�U.�^`�	wJ"TIݾ.��S�!8�C��L`��;���,	��)+	7nc�t�.ø�r��L*eBբ{[�P@4���·��I\�oS��KJ�I������D=�j�ὺ`E�噤���Ϯ��r0N)K�,��H�� ��6M^w`j����u�;�C�-B�1�:��$%��6��� 4Xᵀv����1 �nx&te���v�&6��dbh����;`�Bmo_�
�h�:;�&�#m��RʄҜF5��
��p�ōԫ �lvBȍ���]u�#M\,}����5���l&��P��b<�����,�h�H2?�CLMz�n��gjQ�L��C�13!�l�x�-�\��?1�ԝ(�N>Y��� |y=�G�X#G�+K���7E��@mwW���W��k�0=ٌV���2�H�����~$����:����F5)a�.���h��N�q�?jY}H��s�ǌ����<�'W�:��-�"bM���ӛL�����@��XG|篕P�1���#�8���A�t-�4��(� I'B�݅+"�y�ٿnj7��%K�(��/5�ZN9C��p�����fP�i�Vg����Vg�z�����Y�E �Yh�N
�i�9	jG3�:��c���t�f$~X�h��s�X��HH�m`���C�)u9����ݩ �u�J�*�p�������(��f�`&�bE�$�����צ��4 ����Ci�������*k1W��ӳ�<z�dF�K]'XG$��u����F"���}�@�o�k��V����t���2���h-C{�Q�ω��#��O\D �xUnn�'��
ա7��j� Z��0�qkq�dl�3��ވ�+�ǙU���[0�����V��7��C�,0.41� �]|�d6w�XO-z{U�.2ș�_�����G�jڭ����=q��͡�-*�U��e��P��s6��>��t�:A�Yk�#�^!)x�,l����^&�w���R�eƲ��T�Z0���K����>.�����4i�8?�"�^�ۧ�%egI?z�?s����+�V�r���̤\e�0��,9��n�C�&��x�GZ������V���� ��q D�1Q�R�c�(J�N���R1L�%�y��6�n�nl��"����`yZ��!�pii�"+��Ħ9BiC��L3��5�,@�mm(25k���Wapb���mx|����S3l.