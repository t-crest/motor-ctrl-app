-- DOC_Axis_Periphs_patmos_drive0.vhd

-- Generated using ACDS version 14.0 200 at 2015.08.07.09:58:31

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DOC_Axis_Periphs_patmos_drive0 is
	port (
		clk_adc_clk               : in  std_logic                     := '0';             --          clk_adc.clk
		reset_reset_n             : in  std_logic                     := '0';             --            reset.reset_n
		clk_periph_clk            : in  std_logic                     := '0';             --       clk_periph.clk
		reset_periph_reset_n      : in  std_logic                     := '0';             --     reset_periph.reset_n
		doc_adc_avs_write_n       : in  std_logic                     := '0';             --      doc_adc_avs.write_n
		doc_adc_avs_read_n        : in  std_logic                     := '0';             --                 .read_n
		doc_adc_avs_address       : in  std_logic_vector(3 downto 0)  := (others => '0'); --                 .address
		doc_adc_avs_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --                 .writedata
		doc_adc_avs_readdata      : out std_logic_vector(31 downto 0);                    --                 .readdata
		doc_adc_irq_irq           : out std_logic;                                        --      doc_adc_irq.irq
		doc_pwm_avs_write_n       : in  std_logic                     := '0';             --      doc_pwm_avs.write_n
		doc_pwm_avs_read_n        : in  std_logic                     := '0';             --                 .read_n
		doc_pwm_avs_address       : in  std_logic_vector(3 downto 0)  := (others => '0'); --                 .address
		doc_pwm_avs_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --                 .writedata
		doc_pwm_avs_readdata      : out std_logic_vector(31 downto 0);                    --                 .readdata
		doc_sm_avs_write_n        : in  std_logic                     := '0';             --       doc_sm_avs.write_n
		doc_sm_avs_read_n         : in  std_logic                     := '0';             --                 .read_n
		doc_sm_avs_address        : in  std_logic                     := '0';             --                 .address
		doc_sm_avs_writedata      : in  std_logic_vector(31 downto 0) := (others => '0'); --                 .writedata
		doc_sm_avs_readdata       : out std_logic_vector(31 downto 0);                    --                 .readdata
		doc_adc_pow_avs_write_n   : in  std_logic                     := '0';             --  doc_adc_pow_avs.write_n
		doc_adc_pow_avs_read_n    : in  std_logic                     := '0';             --                 .read_n
		doc_adc_pow_avs_address   : in  std_logic_vector(3 downto 0)  := (others => '0'); --                 .address
		doc_adc_pow_avs_writedata : in  std_logic_vector(31 downto 0) := (others => '0'); --                 .writedata
		doc_adc_pow_avs_readdata  : out std_logic_vector(31 downto 0);                    --                 .readdata
		doc_adc_pow_irq_irq       : out std_logic;                                        --  doc_adc_pow_irq.irq
		doc_pwm_sync_out_export   : out std_logic;                                        -- doc_pwm_sync_out.export
		doc_pwm_sync_in_export    : in  std_logic                     := '0';             --  doc_pwm_sync_in.export
		adc_pow_sync_dat_u        : in  std_logic                     := '0';             --          adc_pow.sync_dat_u
		adc_pow_sync_dat_w        : in  std_logic                     := '0';             --                 .sync_dat_w
		adc_pow_overcurrent       : out std_logic;                                        --                 .overcurrent
		adc_sync_dat_u            : in  std_logic                     := '0';             --              adc.sync_dat_u
		adc_sync_dat_w            : in  std_logic                     := '0';             --                 .sync_dat_w
		adc_overcurrent           : out std_logic;                                        --                 .overcurrent
		pwm_carrier               : out std_logic_vector(15 downto 0);                    --              pwm.carrier
		pwm_carrier_latch         : out std_logic;                                        --                 .carrier_latch
		pwm_encoder_strobe_n      : out std_logic;                                        --                 .encoder_strobe_n
		pwm_u_h                   : out std_logic;                                        --                 .u_h
		pwm_u_l                   : out std_logic;                                        --                 .u_l
		pwm_v_h                   : out std_logic;                                        --                 .v_h
		pwm_v_l                   : out std_logic;                                        --                 .v_l
		pwm_w_h                   : out std_logic;                                        --                 .w_h
		pwm_w_l                   : out std_logic;                                        --                 .w_l
		sm_overcurrent            : in  std_logic                     := '0';             --               sm.overcurrent
		sm_overvoltage            : in  std_logic                     := '0';             --                 .overvoltage
		sm_undervoltage           : in  std_logic                     := '0';             --                 .undervoltage
		sm_chopper                : in  std_logic                     := '0';             --                 .chopper
		sm_dc_link_clk_err        : in  std_logic                     := '0';             --                 .dc_link_clk_err
		sm_igbt_err               : in  std_logic                     := '0';             --                 .igbt_err
		sm_error_out              : out std_logic;                                        --                 .error_out
		sm_overcurrent_latch      : out std_logic;                                        --                 .overcurrent_latch
		sm_overvoltage_latch      : out std_logic;                                        --                 .overvoltage_latch
		sm_undervoltage_latch     : out std_logic;                                        --                 .undervoltage_latch
		sm_dc_link_clk_err_latch  : out std_logic;                                        --                 .dc_link_clk_err_latch
		sm_igbt_err_latch         : out std_logic;                                        --                 .igbt_err_latch
		sm_chopper_latch          : out std_logic;                                        --                 .chopper_latch
		doc_biss_avs_write_n      : in  std_logic                     := '0';             --     doc_biss_avs.write_n
		doc_biss_avs_read_n       : in  std_logic                     := '0';             --                 .read_n
		doc_biss_avs_address      : in  std_logic_vector(5 downto 0)  := (others => '0'); --                 .address
		doc_biss_avs_writedata    : in  std_logic_vector(31 downto 0) := (others => '0'); --                 .writedata
		doc_biss_avs_readdata     : out std_logic_vector(31 downto 0);                    --                 .readdata
		doc_biss_avs_chipselect_n : in  std_logic                     := '0';             --                 .chipselect_n
		doc_biss_coe_ch1_MA       : out std_logic;                                        --         doc_biss.coe_ch1_MA
		doc_biss_coe_ch1_MO       : out std_logic;                                        --                 .coe_ch1_MO
		doc_biss_coe_ch1_SL       : in  std_logic                     := '0';             --                 .coe_ch1_SL
		doc_biss_coe_ch1_EOT      : out std_logic;                                        --                 .coe_ch1_EOT
		doc_biss_get_sens         : in  std_logic                     := '0';             --                 .get_sens
		doc_biss_irq_irq          : out std_logic                                         --     doc_biss_irq.irq
	);
end entity DOC_Axis_Periphs_patmos_drive0;

architecture rtl of DOC_Axis_Periphs_patmos_drive0 is
	component ssg_emb_sd_adc is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			avs_irq       : out std_logic;                                        -- irq
			avs_write_n   : in  std_logic                     := 'X';             -- write_n
			avs_read_n    : in  std_logic                     := 'X';             -- read_n
			avs_address   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avs_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			clk_adc       : in  std_logic                     := 'X';             -- clk
			sync_dat_u    : in  std_logic                     := 'X';             -- export
			sync_dat_w    : in  std_logic                     := 'X';             -- export
			overcurrent   : out std_logic;                                        -- export
			start         : in  std_logic                     := 'X'              -- export
		);
	end component ssg_emb_sd_adc;

	component ssg_emb_pwm is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			avs_write_n      : in  std_logic                     := 'X';             -- write_n
			avs_read_n       : in  std_logic                     := 'X';             -- read_n
			avs_address      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avs_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			carrier          : out std_logic_vector(15 downto 0);                    -- export
			carrier_latch    : out std_logic;                                        -- export
			encoder_strobe_n : out std_logic;                                        -- export
			u_h              : out std_logic;                                        -- export
			u_l              : out std_logic;                                        -- export
			v_h              : out std_logic;                                        -- export
			v_l              : out std_logic;                                        -- export
			w_h              : out std_logic;                                        -- export
			w_l              : out std_logic;                                        -- export
			sync_out         : out std_logic;                                        -- export
			start_adc        : out std_logic;                                        -- export
			sync_in          : in  std_logic                     := 'X';             -- export
			pwm_control      : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- export
		);
	end component ssg_emb_pwm;

	component ssg_emb_dsm is
		generic (
			init        : std_logic_vector(3 downto 0) := "0000";
			prech       : std_logic_vector(3 downto 0) := "0001";
			prer        : std_logic_vector(3 downto 0) := "0010";
			run         : std_logic_vector(3 downto 0) := "0011";
			error       : std_logic_vector(3 downto 0) := "0100";
			pwm_disable : std_logic_vector(3 downto 0) := "0000";
			pwm_enable  : std_logic_vector(3 downto 0) := "0001";
			pwm_lower   : std_logic_vector(3 downto 0) := "0011";
			pwm_both    : std_logic_vector(3 downto 0) := "0111"
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset_n               : in  std_logic                     := 'X';             -- reset_n
			avs_write_n           : in  std_logic                     := 'X';             -- write_n
			avs_read_n            : in  std_logic                     := 'X';             -- read_n
			avs_address           : in  std_logic                     := 'X';             -- address
			avs_writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			overcurrent           : in  std_logic                     := 'X';             -- export
			overvoltage           : in  std_logic                     := 'X';             -- export
			undervoltage          : in  std_logic                     := 'X';             -- export
			chopper               : in  std_logic                     := 'X';             -- export
			dc_link_clk_err       : in  std_logic                     := 'X';             -- export
			igbt_err              : in  std_logic                     := 'X';             -- export
			error_out             : out std_logic;                                        -- export
			overcurrent_latch     : out std_logic;                                        -- export
			overvoltage_latch     : out std_logic;                                        -- export
			undervoltage_latch    : out std_logic;                                        -- export
			dc_link_clk_err_latch : out std_logic;                                        -- export
			igbt_err_latch        : out std_logic;                                        -- export
			chopper_latch         : out std_logic;                                        -- export
			pwm_control           : out std_logic_vector(2 downto 0)                      -- export
		);
	end component ssg_emb_dsm;

	component conduit_splitter is
		generic (
			OUTPUT_NUM : integer := 2
		);
		port (
			conduit_input    : in  std_logic := 'X'; -- export
			conduit_output_0 : out std_logic;        -- export
			conduit_output_1 : out std_logic         -- export
		);
	end component conduit_splitter;

	component mb119y is
		generic (
			Slaves  : integer := 8;
			NumRegs : integer := 64
		);
		port (
			csi_clk_clk         : in  std_logic                     := 'X';             -- clk
			csi_reset_reset_n   : in  std_logic                     := 'X';             -- reset_n
			avs_s1_write_n      : in  std_logic                     := 'X';             -- write_n
			avs_s1_read_n       : in  std_logic                     := 'X';             -- read_n
			avs_s1_address      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			avs_s1_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s1_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s1_chipselect_n : in  std_logic                     := 'X';             -- chipselect_n
			coe_ch1_MA          : out std_logic;                                        -- export
			coe_ch1_MO          : out std_logic;                                        -- export
			coe_ch1_SL          : in  std_logic                     := 'X';             -- export
			coe_ch1_EOT         : out std_logic;                                        -- export
			get_sens            : in  std_logic                     := 'X';             -- export
			ins_irq0_irq        : out std_logic                                         -- irq
		);
	end component mb119y;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal doc_sm_pwm_control_export                  : std_logic_vector(2 downto 0); -- DOC_SM:pwm_control -> DOC_PWM:pwm_control
	signal doc_pwm_start_adc_export                   : std_logic;                    -- DOC_PWM:start_adc -> conduit_splitter_0:conduit_input
	signal conduit_splitter_0_conduit_output_0_export : std_logic;                    -- conduit_splitter_0:conduit_output_0 -> DOC_ADC:start
	signal conduit_splitter_0_conduit_output_1_export : std_logic;                    -- conduit_splitter_0:conduit_output_1 -> DOC_ADC_POW:start
	signal rst_controller_reset_out_reset             : std_logic;                    -- rst_controller:reset_out -> rst_controller_reset_out_reset:in
	signal reset_periph_reset_n_ports_inv             : std_logic;                    -- reset_periph_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv   : std_logic;                    -- rst_controller_reset_out_reset:inv -> [DOC_ADC:reset_n, DOC_ADC_POW:reset_n, DOC_Biss:csi_reset_reset_n, DOC_PWM:reset_n, DOC_SM:reset_n]

begin

	doc_adc : component ssg_emb_sd_adc
		port map (
			clk           => clk_periph_clk,                             --        clock.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,   --        reset.reset_n
			avs_irq       => doc_adc_irq_irq,                            --          irq.irq
			avs_write_n   => doc_adc_avs_write_n,                        -- avalon_slave.write_n
			avs_read_n    => doc_adc_avs_read_n,                         --             .read_n
			avs_address   => doc_adc_avs_address,                        --             .address
			avs_writedata => doc_adc_avs_writedata,                      --             .writedata
			avs_readdata  => doc_adc_avs_readdata,                       --             .readdata
			clk_adc       => clk_adc_clk,                                --    clock_adc.clk
			sync_dat_u    => adc_sync_dat_u,                             --          adc.export
			sync_dat_w    => adc_sync_dat_w,                             --             .export
			overcurrent   => adc_overcurrent,                            --             .export
			start         => conduit_splitter_0_conduit_output_0_export  --        start.export
		);

	doc_pwm : component ssg_emb_pwm
		port map (
			clk              => clk_periph_clk,                           --          clock.clk
			reset_n          => rst_controller_reset_out_reset_ports_inv, --          reset.reset_n
			avs_write_n      => doc_pwm_avs_write_n,                      -- avalon_slave_0.write_n
			avs_read_n       => doc_pwm_avs_read_n,                       --               .read_n
			avs_address      => doc_pwm_avs_address,                      --               .address
			avs_writedata    => doc_pwm_avs_writedata,                    --               .writedata
			avs_readdata     => doc_pwm_avs_readdata,                     --               .readdata
			carrier          => pwm_carrier,                              --            pwm.export
			carrier_latch    => pwm_carrier_latch,                        --               .export
			encoder_strobe_n => pwm_encoder_strobe_n,                     --               .export
			u_h              => pwm_u_h,                                  --               .export
			u_l              => pwm_u_l,                                  --               .export
			v_h              => pwm_v_h,                                  --               .export
			v_l              => pwm_v_l,                                  --               .export
			w_h              => pwm_w_h,                                  --               .export
			w_l              => pwm_w_l,                                  --               .export
			sync_out         => doc_pwm_sync_out_export,                  --       sync_out.export
			start_adc        => doc_pwm_start_adc_export,                 --      start_adc.export
			sync_in          => doc_pwm_sync_in_export,                   --        sync_in.export
			pwm_control      => doc_sm_pwm_control_export                 --    pwm_control.export
		);

	doc_sm : component ssg_emb_dsm
		generic map (
			init        => "0000",
			prech       => "0001",
			prer        => "0010",
			run         => "0011",
			error       => "0100",
			pwm_disable => "0000",
			pwm_enable  => "0001",
			pwm_lower   => "0011",
			pwm_both    => "0111"
		)
		port map (
			clk                   => clk_periph_clk,                           --          clock.clk
			reset_n               => rst_controller_reset_out_reset_ports_inv, --          reset.reset_n
			avs_write_n           => doc_sm_avs_write_n,                       -- avalon_slave_0.write_n
			avs_read_n            => doc_sm_avs_read_n,                        --               .read_n
			avs_address           => doc_sm_avs_address,                       --               .address
			avs_writedata         => doc_sm_avs_writedata,                     --               .writedata
			avs_readdata          => doc_sm_avs_readdata,                      --               .readdata
			overcurrent           => sm_overcurrent,                           --        monitor.export
			overvoltage           => sm_overvoltage,                           --               .export
			undervoltage          => sm_undervoltage,                          --               .export
			chopper               => sm_chopper,                               --               .export
			dc_link_clk_err       => sm_dc_link_clk_err,                       --               .export
			igbt_err              => sm_igbt_err,                              --               .export
			error_out             => sm_error_out,                             --               .export
			overcurrent_latch     => sm_overcurrent_latch,                     --               .export
			overvoltage_latch     => sm_overvoltage_latch,                     --               .export
			undervoltage_latch    => sm_undervoltage_latch,                    --               .export
			dc_link_clk_err_latch => sm_dc_link_clk_err_latch,                 --               .export
			igbt_err_latch        => sm_igbt_err_latch,                        --               .export
			chopper_latch         => sm_chopper_latch,                         --               .export
			pwm_control           => doc_sm_pwm_control_export                 --    pwm_control.export
		);

	doc_adc_pow : component ssg_emb_sd_adc
		port map (
			clk           => clk_periph_clk,                             --        clock.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,   --        reset.reset_n
			avs_irq       => doc_adc_pow_irq_irq,                        --          irq.irq
			avs_write_n   => doc_adc_pow_avs_write_n,                    -- avalon_slave.write_n
			avs_read_n    => doc_adc_pow_avs_read_n,                     --             .read_n
			avs_address   => doc_adc_pow_avs_address,                    --             .address
			avs_writedata => doc_adc_pow_avs_writedata,                  --             .writedata
			avs_readdata  => doc_adc_pow_avs_readdata,                   --             .readdata
			clk_adc       => clk_adc_clk,                                --    clock_adc.clk
			sync_dat_u    => adc_pow_sync_dat_u,                         --          adc.export
			sync_dat_w    => adc_pow_sync_dat_w,                         --             .export
			overcurrent   => adc_pow_overcurrent,                        --             .export
			start         => conduit_splitter_0_conduit_output_1_export  --        start.export
		);

	conduit_splitter_0 : component conduit_splitter
		generic map (
			OUTPUT_NUM => 2
		)
		port map (
			conduit_input    => doc_pwm_start_adc_export,                   --    conduit_input.export
			conduit_output_0 => conduit_splitter_0_conduit_output_0_export, -- conduit_output_0.export
			conduit_output_1 => conduit_splitter_0_conduit_output_1_export  -- conduit_output_1.export
		);

	doc_biss : component mb119y
		generic map (
			Slaves  => 1,
			NumRegs => 8
		)
		port map (
			csi_clk_clk         => clk_periph_clk,                           --      clk.clk
			csi_reset_reset_n   => rst_controller_reset_out_reset_ports_inv, --    reset.reset_n
			avs_s1_write_n      => doc_biss_avs_write_n,                     --       s1.write_n
			avs_s1_read_n       => doc_biss_avs_read_n,                      --         .read_n
			avs_s1_address      => doc_biss_avs_address,                     --         .address
			avs_s1_writedata    => doc_biss_avs_writedata,                   --         .writedata
			avs_s1_readdata     => doc_biss_avs_readdata,                    --         .readdata
			avs_s1_chipselect_n => doc_biss_avs_chipselect_n,                --         .chipselect_n
			coe_ch1_MA          => doc_biss_coe_ch1_MA,                      -- external.export
			coe_ch1_MO          => doc_biss_coe_ch1_MO,                      --         .export
			coe_ch1_SL          => doc_biss_coe_ch1_SL,                      --         .export
			coe_ch1_EOT         => doc_biss_coe_ch1_EOT,                     --         .export
			get_sens            => doc_biss_get_sens,                        --         .export
			ins_irq0_irq        => doc_biss_irq_irq                          --     irq0.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_periph_reset_n_ports_inv, -- reset_in0.reset
			clk            => clk_periph_clk,                 --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_periph_reset_n_ports_inv <= not reset_periph_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of DOC_Axis_Periphs_patmos_drive0
