��/  �ϭaK��9#|1�
�U��W�G?W.=EE���{���U�#+I�X��aF!����85˒���TDW�R�<��^�	ύ4Xi�&R����8U�j����/|� s�^�v䅀8�x^�
��S�Zgw�Q�	[��X��w�h]�ص�ޙ�6;�6���(��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[�Ţϝ�(��N���b��Pe-�-qE��jV�$���e��S��/jk6N5�)�y���pA*�H|Y�7P D��|JD��S����"c��&E���\�2������Z�uT�x*��%�KaK��;aO~E�5�Ћ���0?��%��	�.mo���<���̓���'�J�����6��Y|���)C�r�,������^B�8'uݩ��J������#�kg����QB��m���dX7��	w��V�{���H��a�q힖Jd�h8�р�}ײ��w�'��+��Ta�!�P�J(Cy:�Fx�ߗ�p��^�����qjԉII�8�$b���33���#	РO:�*��t'��-��	�X6���O���8b�[�W'{�8�Z�$r(�Ρ��<��#3-q�u�5T���*ez���d��7��ĖԄ0���p�v�O�-)7��.�?q�h�FN���,??������z�*���P��1��sb.I�z�,�1y�)�T�k���u�+u[���J���1�r�M�hhM�Qs����`��iW,�����8	���g��l�,�{�W:8��0��"`�vE}oY��2pJ|z��M'��UD�m���oj/���|����))����F�u����.��g��ҕ�XŽ&m[;�1�4L��A���[��tX*Nv
�q`���8[���l�?�g�W��G=�%cX������95�󩰖e+�[xK>Jj�c�_��X�d�r�~��G��Pاmύh���\ ֪q:	�s4z�:�*u���
�`�#'�I������)��q�D $�Z����b�K�8M��\>�)�2�U>ݨ'��K�Im��~��]�6)�B�J�~%�F��r{�a�t ��m?-��%�9�ݒV�_�ŪAF]�����<�ʺ�-]�hp��UD���w&�g��a��Y;�X�2^>�҅�F���j��s��U��HeU506�]P�=���|p��N�&v���eQ[&b��]�����=.�"jsg����AӲ2��cbZ��Zg��\���ϡ���60L��v ��2"3T�SXF()�=�a��|!�8ʴF:ц'�W'כ:���6o��4r�*i�Y�"o%���j'�Ta7	:�Bѝ�����e��C��8�M �^�9f���<��Wb g���ps��G�$����}�S����3�mcKUz�����;e�}tlSݯA��\�ք=Z}ݚ^���*p�6����-i��cOB�����ƚ���$�`�}��w�2=�#\���f��z��ъ�@sUU�9}8v�o���R�P��ijP��Ǟᝓ��[Tl����\��\��X��R�#{n5�W6?��]
�$�iĘ�9���b�wpS�טn�G��b�DN�|U����j �1[���"�&b+��A��r�`�!	�@HaSC���eDg��)�6IJ�rP�W������Dݜ6d���c��@|#}v݌�)n ��,N�2S�S���P���ܕ�A�2Qil�%�)=�~�C��|7��&��]5�I�쓺؈�Y4�m�nG�M�ur%.�{����� �N�������A ��MYT�}݁���-V��ɥ���0������	�L��u�Hș��e+�����9��*O�}C�E_�s@�6թ�r��Ά� y4h�_�\�߬p�sk��J���I�`H�s�C�գ��5���m��g%�ၠ��>zL~'C��:/����F�`Nr{��d;�J���N"�%�
�S7s�9���AU����~������Qg�����}�Qp�Ä��%A�{��Z(O�o%u �8��Ƒx��{e�q��X\v���tZI5� M�u{����܄��=eq���~ߟ�1��\��;����љ�]��������5�]�ά X��e�B�B����7Q��9��I�q`���}KM��FR����a�c�k����fGQ�t0����/�]��(����$o�Pg"�T*���!ib�`JQ"br�0�E�&�J�KW�ć�=��TL[�IG�t�}��u��aoX��h7�R{R����=`]�B�*�����h��m�W��Q��2�짆�an.&t��sc��ߔ��+Y�4�fX��t+��Er���9~��k�7ϔ
Xр�]~n�9K���t����`2[V��ά�Mj���H]�#����d b���S�P�йݏ��p�����Y���@~�:Ԕ$j��5(�BQ�l7�zT{?8-�q4����2�.6��p���JqDU��s�m�r��1I��<`��G��DXt81��q����.f�M�8�U��@"'4��3Oy!�*�g��(g�	�l4/X�qr������D���*Q�5�T�;GI���V�ԛ/�~T�U�2�|/Q�x�[����v� 6�������/�0��s
���)OAca�%g��C�a��Gub��(i�s�:�yU�w�iJ��8����������3�yv�H��듕_�KC86��1Y��g �b�V�<�Wq��-�L&����&������w��|."%�y�r�i�0:r�6��{"�J0���-0o �َK����6�����Ӏt�HY>$Jۏnm.�����U�M@�m��-��8�ڄ/{ϕ <���R�Z��L�0!͸5��m-�of��ɯ{x2���j+
��k��;^mD�����h.h�K������ax��*��'�\���'#�
w��}m+ӹ�?��/2�Tb�q�\uA��nWY�9s�9���I�dQ_�`�����`���<-w�h?�6Z)�h}9@5RJ�2�t��~��o�w�M���qY
���"ʢ�т϶�ܸ?�8N��-Nn�d,�v	��Zd���M5��H�Y�wfAD��#x�����8�����9(6��6+�����r_��N.v��KX%���沧b<_���K�2�P� w�{�s��e��ިk��s�h�w���b�-:���˵!ۃ��1�A������#2P���0l�]��ec���B/2��
O��+��ջu��	��S���g��?���X�"nh֎�� Nȶ�8;p��cA6;ӄP�P�Y�}}V�q�X���*E4?;^�«Ő���4Y��
��:ፀ�����s���nz-A�؁�.sy�ĕ�-d���1ଷ�->�W|��xj(c�A���L�.3�}Lm�}$�o�2Ɉ9�Ep	�A<z:���TPkbUS�:$3�]�P��P�r(Y���w��z.�y ��X��_t��������EÑ]d��ˇ<䤔8�Nك2)�;��X�EV��ܗ	����C���B� a�,��(�w>3�K�=�w% ��)^"��B�Wz�
��Q�9)w}3��������<Ъ�ņ�Э�F~�[�z:V�%xk��ʻ�/�����c��Ȼ�ɍG�0�7�+�� A3/�P��ƒe��A�wep���6�����H��rwm�����j_���{m�*��q���ݝ�)�#���j-���L.�c^�/u�S���43T�O��d������}
p�u�!|����7㋩�]�gT�ʇ���tJ~Ũ��?|�n�7�Q��t�ג�� ;gwh�u��l�Қc�!QO�I�f$� �(>ʸ\�u��.��4��ήIl\��,���,�?k.�/���K�3pk�q�*$�gs���'
�r^XO����y\�'d��X�J�@�a�R������8=
�O�u����7�{�Ծ�2�.%[���0:W�S��dεM���cM��0� �'4��z�������;E��j��x����S�'Fbd va[�.p���
1���]�������_w��
}lg��#�Hm�b��盕$E�Q��p�����eAa?�7� �9�'�7 ��2K� ۰����*w����"-�����Ap�Џt 7��^r���@������&�Cܼ��ȕ�_y�
�%����g�J�w����w�ghߧ����^��6D�W��eDH�
��&�@I�=B?�+�J:���.��ʅ<#�7D�)˝C���n񢟚^Aq�95S�w�]"�*��D����4��i�__1x�~�2���k���60zoƅY�5r��b�|�c��S���b�+W��&���K���\Ѵ�k����0"z>�f���S����������N=��4D����گ�1U�߽�"˸>�_�`ea'�,�7��ǶM��N�c� ߐ"I��T>�T�|�J�c*�*O:�1�OW5O^�Kf�4��Mm�O)��P�٠$�zr�U}�w��ٚ�L{2A�͟����1��@Z�,hc��x^�®���L�]8��!,h&9�闼���u ο�����K3���ڷ���lQ_�j|LߦeI[����[��{~���u�*��F��{v��:`$���3Ą} �6	���3���C�c���:I�����wqA��46]iu�a���0�5�Xq�n������o��t��ǟ����^U�1�D���H8ԝ��_	��x����6��{,V����+��}X���9�I��l襯a��_Y��b,�4��#�L�?7��a|O4y����Ӂ�e�G�1��16O
d�d|���5�ȭ_�-�BK}��x����/�z��ɩ�}�x�|X�{yփn�N�3<�ty��̒��c�.����\W�#�Ma�|��v
��l-*R�	[ ̳pF�8C\�.: )�IY3��e:�;��㫎�WK�N�|o�ͮs���s�4�柟���~Jb���*���[��
�_��5В�1R�����?��*��N�����m���	����>zDHL%"�d@�m�e�OW�!('?��,r���K����=����<F2`Zm+����B�(jƄ�:�Vl���^˖U�Tӆ���fŹ$N�3;���ܥ��,:J���m����^�H����ȝ���)�`��36Ea��!~qo���-RY+E�����gF���&�h��_"�eY�(�d~OS0q�y���}�q�d�z��q6�!�i��M
�41�$�>
��\�����ڃ�?��+�%��W����Q�#�sg7]�K��5^u�w�{��e;� ��vY�"�<�hA�ڬk�l$4�,!�AIڜ��2�\�Ҝ�6�ܼ��@+��$�>@�ު��C��a[��&0x�!�Q���[��Ӻc0�eXd���	�"�&2h�vn���~��� \�=��bzIg�/��2K�7��u��ҵÓ�����R���$ۋf��%��r��a��K'������ �X�X1i\���^0R���[�GY�]HR����T_��������~7~� ?&kr�Ꜵ!�1pVJf3j,�h�j�,�"���gE�Ӓ���u��u���_�%�\�1D�e����!k������e�<�l����
R�e���	��>�X��]�ؤ��a	ch��S-�<R��:�uY�1
�;.������B�@S��!-���Ԝ�^Ӈqf/�^\��y�N��,���|�7T�:��/�S����b��̕��`=�����d¥2$�~ �tj��*�wѵc�>�����C��]�:ki�N�NL��{A�5�|��6�����1�=��� ]^8���6O�0W�l��<��y}e%�Θ `GtJ�[�<x�RS���6��QE���
�ų�<"?��Z�>r-��C������Qg��;xFo�駧�wWTj�;��j���۷���)��^�憀�u�����2�T���_t���HnR�,������۴�=(?j�����Ƅ_�ѓ�]?CL.�ΦuJg;�@Tp$����'���?�˪���
;��.�ç]�����F[4�β-X��~�ۨ�T�SUu���}��C��S�?0�pg=�8��N~���o������o�A;dI~�� ��瀕yE4n�AG���Ƣ���fK����B���f�ܣD��+�W85%��t��T�Fn�����5��ţ�$1s�(�`�rmYg������m��v7���Y�7�
��n���`��e�!@̤��5���O�P��<�~��ӱg�U����d=�T���LM�)��D�<���`t���2��D��������͛G�B��^i��^� ����a��2���t%�3��!��v�`$�c�L�O4.��/QY�<��z.�AZ��a�%Uo!p�7���,�i�:�W��M4����]*��U`��jc��4ҽg���^=�o:GH;�zW�e.�K��1�;R�%�W\�G��(he�S����~��Vt$�h������:�_� ᬭkuw�(�l�u+WǄ����A���l�W,���RDc-`�@�vL��3����j/p�
|��NU(t��d� �~Q����J��l����߬�lOmAjɟt�cӼr��@1�R��j�?`��g�Y����O�2�9����y.3�>�-�6bV��+���c�đmx�JC��i�X�9���2/�ӡv��-�x73�O�
vGҳ/^47��-���U0�E1l�^��gBu���C5xc(�"��>�Bɾ�G#"�Z�o,�z���ۏ9n�Z�7h�FЍƓ41�m��AE&I�����]���9���SpG��ʴ�:�������n仔��o0!+� ��nt.꬙�:	� kk�VT
<�,V�K��k]���I�R�[�����=x�%@�r�̘z��?w��&2�S���c��ņX���""�d���ڧ8y�%e~TъUR�mX$��F�w� V|�uQ�����5���/.�a�"��O���yi�k�e陬�SFV��>����2%k��6�i�|�0�w�u�P�^2�ZI�
´��qwy��>{�;����
�{!�1�Ŀ;C4q�u�(�^�q��FcO�R���Z�o�Z╗��T�Č��ǑONLx�K�p]���M8�����Z�q�:�1ґ�ZgnV��bB|�A�m%\B�x���IʨȃF��}_R�lйt��8�y���
�+y�ݺ��ڳ���}�I�b#���%������J�������ƨ@`H 7QBH��Ԫ��v���k4c��#�,����~�-�õ�O���x��g��~��</	5��k��4�J����O���ì�k�e�}^����1���E�f;T�0��j���*��W�S�A�&:e���T��}�bňr�����;C���>{NQuB�.��[��r�ㄍ�5E)R3���xJl��.�U�m:xt�Y��X�f��;��>:}
+�]������Vy6W�!�a��'/]����>u2�h@a�a��11�-�#�j��E�/9t��S	洩)�.@���]�0�T����:%"ݡ�k[�NZu1�ip��[F�4��C[�,��P�y	�sB���ls����0fX��L�
���%|ˮ����l[�0�5�h��*)����eޠX�_��&�q18c��I�Q'��6i��VT5���DF���'3Թ2y*�'����۫ͽL�χ�����6��+��!=�W�i�!T�]�Z��\�]~#�R c۩Npb�+u�̞b ��2&\KIq��;[��{BOnk��:c���r,7���~�U
Z�!����A�jc��\2��@:���E��t��AM�l�Z������S��>{�&ul����4-fw=e�"ڤ�x��}���w9H��[7F_���Ȁm:T�*N�O�G�]?kp+��u�>`����ɨp��w�1���)#M"x�NܝĚ��Q%�i����*	��c�fo��1���Qg�<�9�� ��������vԹ{.��έ^PW��]�TWU���3f��%s���U�̙f����Qf�e���;Z��к0�"7���R����w��R���{%#ӂ�s�ѧ�=b4���oD�B�6��j������f/�(dW7d��z��'KSB��f�zǪ5`'����T-#�kX��|#����Y�l*��Cp�1�k��!s,:�#i�
�ԇ�&zMۿ�Uhw%�t|�Qz}\��x�ǲg�c��V��t����#R��\�T0���l�aވ!S
�M�p<�z�^�:���X�:�tc�g��+�I;*׊R���a�wRsp���>�u��p��il1��{���,p�F> ?,�	���*��FE��qp����2˳k��Y�����˻�N��nm!�ߊ4<C	t�6TA�����a�����?hy<A��?���X�����ʯ���aݴ��"yV�7�+��}&&'�`ʝ"~�Dr�|�"u*UZ����ߠ�n�	21�<̊$:�w.�w&�������t����Sm��$�!���l���N2���HTA[3�.����{R�]�fj"^6n���sMɭ*�jL ��ˤP��=��v��$�vyǋw�6*c�mv������]5��HF�9�B-m��8;0b~��>u�Ф��T��i���`@\��x��*�:t����z�L�˔|h~�1�fhVا� �Z(�0{������(u�3���ﱷ+���k9l����v�|J�d`��ŵB�	]*
s8���i^�'[ .8�Iù����M���XX8D�3_�zd���M�W��>2�7 !F<F�:�CX})�+��ː�D����1y:�N��V%�mzf��ﴊJ9 `P��>PW�i�ػ����>Y&_@-ʽ�/�]DY�zD{�:���鏽�k�r�ԍvN��$5P[��q����� ���P��-�׎�F/���j]44G�^���r/���� !�v߰tn���m��⺢��]>X���������vm鴀<,��Z���!��F#b�-�C}c��R�o���j����z׆w}7�YT��[�p��%���ۋ�����ojn�Lu��7	}&��溋�)�t�^�;�ݦ}��&)Xj!�ǐUӋM�50�v5���$���u�O�\b�N����̆�i]6�09}ݷB���_ە�N"�	����<��9�3��a�	��.���Gu��SǲGU�+v�Y���6
�a���C���\=�w�ǩ[{e��
��a+�6�1���q{\<�[
$E�L����[ Q���2y'w$3{	&����umwӂ.�Ƞ�,L{;3Y���ci�����4�崌_�;�S�"���,6��������F��0��U�i���Eq
)���6hG$�*j�.-�9w��ɸ׈�	�d�y���+��ֶ�1����k��vQBB���y�|�[��uƔ��eۏT�6�ý�O�l��X?���]\;r;���x�!��f#B��I�m��+�˔��c��Ȃ�Q���j�E�bJ�vm�� ${��'���P��ɳ�q_�P&Sh[��_օ]�KJ^x��EY�����~&��(��$:�x�9X��h��L	$e��e�o�(1�+<b�|����Ϸw:��(n���P�3# ��o��;b��%{��	w�ikja�H՜��G���ᮅ�y%oH�=y��;���'�W3�{��W��v/Z��$�:���u?g���INX`@M��
�.{Z��n�F��7�:l��~8
����t��%v� !GG��j��ois[��<ƾ�i0�5p(iw��z*�Y�SYm�uW�E%M��Vrd5`>��6�$Mw_�4Vӻ�o�����Z!�Qu��Ti�P'1�߬��0�Z�^�A�lލ:�EVJ�\�>s�9��k�P�Ӌ���?�jY���>�;B��.��!
h�p�~�OR�7���6��o���t�	M��>�i��m��I������
�A ��s*�żz���/i�Ɔ���ZY�^i?��a���@+�ָ�J�qQ�T�)3�䜻V���v��6yy9]�~oU�	 ���D�E���y!�NL,羋����d"3S63Jո�s�4.�#�U�vDo�v8�Ҭ���#��C�Zؒ�����Ud��B�Q$mu�I�����j4G�*�wf>f�ڇs��WnN-��ԕ��a���o��]� ���Kj���r��������p럎���vY_d��rϯ�����H�eOZQ?�[�JՂ��,w����]1
�¾�d�ֺ��{�(��ZL���hv���V�<Rbw޶]!��9w[$�"�ܼ��o�����[�c�Y����}��H�W����`�KN��wQ�P���}��+O�̎�Lݔ���!ʛw�BZ����j,��4�UN)���u$1S�O�N���9�!��l����:��_}͎�-�io4��a8̽��sL7(ƙ��n���'um���a\��6����߼7�7����kb�����|S7ؕ���/�B�A�K��u�ѳT��0*����̾g�l:�AWJl#ٛPF�R)����'�2
��pM3nm�<�*�A\�IK!MUnԢ�t�j�����q�U�hy���.T��cڀ������P
��.��O�l��3�M����a؉�ivx���0{�jk�=3�b����#k��g�����;��s�F��--D������T����� w�'�*�*{���3�����$��a�'n$�ū�M5ҬV{?/�.3���@�RNB+=Q&4c�+T�`�ƕ�z�{HS�Ɨ�Ԡ�۠�h��m_F������/��a��� ���S�"��ߘ�����Uiu8G�M:]kH��WޕM'ǭ����C,}����u�;�}�����! �œMhŪ��S���bپ43>�%��m��н�wN�,F���>�6�X{(��
�w��L��ѽ,U`����ni�)�����1�� �\���R�nB�.�h�� �$gYZ7��e5��!FL������e2��ni�y!������U��\��!�R �[r(4D9GWC����WgȠ�������#J�/��O���|Ɔ��(��V_��ۻ���}yc��|I����)��W��8�7��V̎�l��QK[��[�ч3YS.�y���q�v��yà�
����5�ԁ��ٌ�h�ڝPQ8�]�<�]y�:��� `5�f�-h�a]�ͤ��K0�>����oNP���>E��Ά� F;�vQ�
3��k���.6e�o+��a��}�k����N��E��6�)p�Pk�]1\?3sU�ݓ��ub㒼ABuBv||۰&��$�f�U��6ܱ�6���������Ak�L)��Q�y�n�+�O��T�XL}Z����:B���Lh��*��b��������h|U0D4V��3FO��y�R!��륐2t��!anh�4�B�M���jf	����}̻QT�V�b\�i�Gӵ�'t竷�m�p��ڐ6Ro�5s@TD�~�(��\j����6A�M��Z�i��c�	�;j>���d�E\�r=�I�;�l���mR�VEk(.�P},-�}_A��$�
�0z���=��4U�c��x�E�/x!�|�`��^R]yS؉K�!�	D������6����aގn��KZ�zE^׷?&�Q�?!L�`)�Nt>S�K���Vt���|l����	ܯ</��"}"�֟�+����N4=��":GnZ���x�GD�^
�[�>�p �k����P��@��I�>�sI�N�w�]}5!o��{��/�U�:�E�2���ɐ�7&	8��3sŻ��D�im���k�1�u�V���=!0UkZН8�}��b�@B���i���F+��Ux6
ܾ��XC��G#�)�~Y�f�/�[_n�~�SJ�A���Q�T���1G�gh���8�L����&��w�-�>��J�k���+){��+�^��7�R[��Q��(H􁧶	ʑ�7���4�{���v�<&[C��ߗTɯ��a8���|����y�M?�feܔ�a�#�����:M7{�XG7n���:W�-<��ʊ��OjzLt���ܞ)�o3}�����-�þ�n"�m�(0��N �O쓩�fb���!I����J#�l��G�����PW��I�h�wd�ű�(��	�ڠ��Fg��.F�V�N�n��ecq��a��F�;6b�Sj3��"�)��jF7��~�<jʢ��6�|l�"����.�"��A3)�\oO
��1�	�+�̲���.:�ʴ�z�]�$�MA �� �{����{F%I�P[�E��V�u ����[�#�x����
�t���DɹT��>�n?w�aY$���yY��Lzbq씰���է����I9��n��1�%ѐ}>���@T\���n\����{����h�&�r\̌
:�z#� � ��K��~X�#�x�PT�P�U�Z7Slz��QM�e闞�r������
z��#3jL���3k��\l�)]7ÅW�I=�/%���ě����=3�>'��� ���ם��?Ro���x�y�����,�%@��	���؋j��!DZ�J�P������1ƿ�ck���@����j��,w}&�B�A�=�_O��:��f���=��[J������b�
����C��0�\D�"1w����Q��y�i�.�xbIJ�QE{�e}��.}RՀ��)�>D���B���&�?���g��c8L�~�(�x�9�d���L�V;'�![�I��r��)�6�ֆV4�E�4�H���K���ᑿk:ň�afX�y��o���Oغ1��i�j�����tܦ�Tw�*5>��:�%oI�%Z��E��c��< ϛ3~W`�GBh�ٛx��m��Q';^�{�!��v����;��S����x��j�I����#c>M��y���膜�l6��HI{W�g|��E�KX���5�IQ}���gk=Z�~^5xQ3�����1�Lm݆9�f�8	Pr�ȹ{|���/Fn��j���E�ێH��_p�-g���JbXDb�TUT��4�u��s'�nש���懯a�s��`+����C���C����e��/�i�8u>0���>��Wt�@�Y�$'�x�ML�`hr��w�Ǿx�^�<Y�܂ٿE������E�9���ή�-�)�d~t4�] q�1_�
X��(�%;��V#6�=����׭j� ,�����&���p�|BL:��D�-��g�[U�.Mȁ�����3[Q���xEj��{5;�W��vº�����Y����0j/�7��H��M{���Ȱ	�hkYk����\���TR������1��[`%TU�'�)��
�B��w�wɈ�;�.���^w��0Wc9�\ہ &�4�I�*$v'�
~?��a�p���'D�-��nIA�sXr��ؚ�&<���p<�P���쳐z��.
o���L�xq\���43��u^vK՟��S�6�X�9��o�Ak�|f�F����Be���;9x��{=�!�}���@�	ΰo�_;b��evX�Q�%����ohF�En�O�| ���P��}�r���5��n���0�=~�t/�F����y��Oo"���2��ˠ/��4�Y͖{�ӻ���jH�⡉�q�c;��a�[
a}������V���x�R�P@����\z��(��An r��ݏ,�����K����s�e O���z+���o����^��Q㠣.��\#�4�Ѯ��4G�]ܰ���s7A�ʎa�]�]�W��KE$����{uf���V<����&{J�ڌ��7��XC���ĭ�CL)���,dh�Tڰ�j���M���\Z�����GuJ�9 �#��*�֎d'�Mv|QG��r�U�::X�q�KD<�nz�S������������.�yܵvC��5x�G�ysw��j�.~G�$�y�}x���<]�<��%�*����3�V�ΑF�i�u󍨐~ o�u�Mh/^��d(����Yˆ(��X�=�b�܊�J�.!�ʤI0���r^;�ta鹔2x�8m��+5���M��U+����&>Gi[���t[w�`2�A#	>5Gn�KL��Y�*�N��e�f��!do;R��B]!yXǹJ�d��m2�Xʰ���_J�S����È��<��#e�����˝t VĀ�8K���> �����gyb�BǗ��RW��P�׿�O�Y}�nI��8�%>�ɺ�s_$KV)cr�ٮ��?�-��05c�B |���X�F|��?>�~�{8��8�E�e���~ݒ���IA����^cb	��G�f�+�pYƪ�K<�.��i������=u�b�w��&S�#.>%J��ڈ�8u��/�p3�dySNY��Ā$���偝�.�X)�!���j
{�ś�}]^��֧@P���@^�G�$e0,�����(�i��ш�*O	��w�7�yyE�����^3MN�}��LO=~:u,�ׄS��ρ�D��i�)���۰3:�5Kd�jw�e��7i%��0����<b�2�OB�8bR|@P��e�G\z�������V��4�E�f�M����84���Vro/32H�k'{g�W���*)FD��#,��r������x�ѯQ[�4�'Ėٌ��))�A
��2����e��4�zkv�rgm����� jO=te��32�M�!���Ȱ�g��Ez�;�M��K�xA<%�(sg
W�`�oe"�2��r)I�'��R��������Wkq���m�*�A�9�<:��J�P=����	*���4����ͤ�!�@��]���U�.��m�\�d���!��s��	�yP]<�Lԗъ��(A*ӎ�Q���>�	SlT�ͬ5޷����.B�ca���g�2��hEj�kw�O�q:ք��]o0ƺ��q�2q�!�)���LH���[���m���|��:�$P!Ej%��0"���5J�B�Xe_ �4{L��V���kRO��-�T��y�X�����D�j�C΢f(Qd�q�����&�;��8��v��%qf�ܿ��zq�\`7���'-'���o���WîRe�%E�`�&���)�x�|��M�z�ϳs~�&�&�k���[��w^�
�F������_�K6�$}��r7��ƞ9�s]'	S���;A�m�sNĻeGR�`��Ѱ�������$Z�pJ[��#:)D���� �E���w��{�'���҃v�}���ߛ6��{�B��r|��2i�SU|��1�&t��̕0L*�8�TX�2��#�����h����gȔ��Gafm�bGț]I��+��+��ԏ�X����#g�地ώ0V
���st����+!�����ӧ#1ves��cB,��/��m:�F��ǯ�p�@	��e�KL����_֫�@"k�>�5��!b�Ф��xL�n���cħ�.����8y9��ݎ��f� ��*�/4�46+T�X�(���z�]�g�0���3A�[�\��lˊ�����:��c�ݟۚ5�gg���c��％bm�����Q���n#zm[�x']mo��� 	�:,���=����n,����LZ'�������MM TB��Uyڢ�氼oIqd�b~[4�%�]Q"C1��`��uWi�Oq6�`�Ʋ����:��c"�c����`��Q����� e�)�t��"���� ��aX�n��J��
���-�U;�ȴ�h�.�]Ħ��g��N�`�4��eQ���,aW 2�	A�Y�i�0Y����ZvU��,���^�ކ�m�$���@}�;c�&@ȡwe�9��`ɩloGs	�jQ���v9���[G ��ӌ0����^V��ۖ&�f��;�{"VCP�A��(�p�����h�8�;,��a�L�r����º�~��)"-I.���*<A6%��1�9��<�J�V_6�BX�Z�������*9�N��V�f�:�J����k1�5�H��$!&���cK��$}S����J� h�\Pڂ���̉iF�}��ԷF�	��d��}U�CV�k�Mt=�V~�RrY���̍1c!�4�ڒ5,!Xf~P���f��z��3�N�Q�d���FG�[�zH����K�b�����|�J"_Ç"��T�x~ꉬ|��&rf�}q%u�c;�{��[2�Ә>7_Q���>i����7�ؔ�xٓ��3Q�0 �����4�um�vfQ����U���;�nY7W�)rV�퓹8N�n���g�D���Vw��Jp�7�K��#�-Sq�' ����>�y�$�+�S�
��S��K^��ĵps��6ow\������<�;@�穀1�S�8�FÊU� ��줡��	װϸi�-� XM*`i�� �P���1l��P=���Sԓo��97s�7�WJ��t/`�>x���q1u\b2i��,F0�]W�,Qt}˘CԌ���)��-�
̸�+jq\�h�Z�1`��Y���,���}p	}Z`b]����U�
�X:d4�Q�+���a0�N�T�=��N�<�-,�E	�͒�Ꜽ��w[�7Tpt0)���.�Q����֨�U�e�3
���o��h����V�.h�����Ź�{.����W8�OU���^�s��9
+Bf[�O�D̟�K�	|ͮ�X^���=HW�r_�V.�2�Zn:R���S��Ѿ�̋�o��a�u�ȤIGNe+���bL������6�djA��8�I�f�M���ū6�	�b���@����ݝA^�tW�F��:wU6j�U�zoP\)IP�8��a�UPCt%[i�i��6����%n��}�m��[��)*�zE�d-![�)����x+�J�j�&y1E�bi�)���s��4hA\��r
�+��H؜�<�'��\��aPO9���� L����>��p�39��6\�m�4�	�/Z9R᷁l�B֑��J���I�.�(�cw' ��V�4���$����
�u��W-兊l�\A~���G]n���p�f�?-�nIw,�dY��9��2FQ-5�/�ИHy]c��<ߜD8�;���6d��-�c��֐8�+u��	�)|�)��G5�$��׌j�t�;�#8(����qEŠ���F����x�ٝ�C��V��m�\_M��(�V!xn$�9��9���Iɝ�i�,��k��/��9��� '�d|~�:��ؕ);
�&�E�������%	J$�|Щ@l*�T.��>���W$��1�hf��េ1�D?�����m+�:��ب<Ss�ε��d��F
��1�yF���K��6�.|���}��R���o�F^R0�P��9ȗ	��؋�����XTڻ=��e�䪵-�U���R�J�o\� ��i���gg�h���
�P���� ���)�- �0�t���=x���<�f� �s;5oY2�Q�%�����C��,!��L>!m
d���)�{v�JЮ�'3���#o{�S}����?��D�JA�?֞��'O��y_gʠ-���KH�y���ΰ�79ȟ'�8L4��Q���O�EpãOVN8DI�Gj��*��&e`r�wxF�!'ͻ2I�{l��pT��T��[�0ͦ���J�� 
�c�_�}|��z`΄�'�?����ڝO��C�.�Xq��ՉO���p�����#T�����we�R�)���
�v
$�!L�q&��H�Ӽ���B��mnĉ^���̘v,��\��;�E*������p;:�O}.lV�
o|$����{�3S�5�ݖ?DD�#<L��Ё�V�A-���\�m+)���uP���������"�*������t%�+خ�7*c݅�T��j����7=|�(��@��R���bfvй+|H�m6��'�$Ɇ�L������c:��Ld�N{�� ��Z���z����#�K�D�n�����=�<��?Y����k�J�����AcOǱ������;�X�Y��˰���Q�!L����ژ�7��52�mޗ?��4vTS�8��?��w࡮Q1�XR�`����\�*��b��u�z�e���ʟXAD��d1s��a�s7l=ϧ4��q�l�O_ļ�-⣤�26�Yi`�N�k4���^�Z�7HGŝrqs8��3u�2[Z�z;���!�z*~T�'9\@��Q�+�%�����<@C��(�F�ȭź�V}f��Y��p���fLS*��/絪5'M�S���Ĥ�zW.h[U��N���%dBL�N_�ٕ��a#�Q���GŤc��3q��q�d {�>L�펎�_�u�n[.i�^�"q�r �b+��9Qy�vWq�ɺX�=���F�kX6�)+�d�J�Ûk�hRV����"�k�s�2ZdC�Al3	 �xxgu$�5��E	�c���U�X��#m܅_u3¿�g����I�vN(�A[eK\��V�$�2{��t�Z$� ��e*�QH�C�LZ��0vΝ�1�l�_j��� 7Ex裘|��P����$��`�$�9E�>^s�i�7❯b����P���d���}(*��FYU6��N�X�F�lƪ柒���to����?��*����ڗ�����zE0}W���%np�b�Wisr��]R1�DDm0R�n9�N�4ٕ�/��ǭ���͔�p�il�U"��r ����)uz��NZ������O/`����6�? ��]x�)Oō���if��\�EFxaq�2!��@*�s`��<˔q�oY��n�>t��򩰐��A�J =I؏F��1��8��(*�g�b��Tr�?���!V.`
�?�Z�� ��E�{%IB� �2���!�:$�zY*nŹ*�Wp �َ��ߗhuN&\���j���L8��,��`�$
u ��Bχ��vV�9n/��&	���Ā]�5Fۗ�������X ������e5����"au����*���ٍ��g���&�m$�n0��	 z�浔�����Zg�̣��"q+��\�8U*�\�C<��?7��A�!t�@����Fg�R�B�mY�)ފ�,�nX����D@�*�'�˷�9�zo��#�$af�?�.��7�W�5O����U��������w�wt�u�28G�\� ����܆t� �؃��ʸ�)|�o����*k�TAK�i�y���+�CN�6He�e�\�;�����:��=��VXl�V����g��a����No��5�rG������Y��d�?�E���0�K�Wo�/��sh~CEִE���Pd��=r�+n�Ϊ� ��/����>�����{�5�,�L��$�#n��D 0Q��}7�����JJL�r�T2����/����8��Q�R�'�w�`�-
@Y��wx�=���_�y��#/�,�wxU�b�#V�e�G�v�X��4��EQ <���4�Ē�dطV�i�i;��N*�-��p�p��}��WI��,���fG�Έ��5d�A�^4�Tgz�Qf�?s�y� ���s[:J�g̪M_vw�j��l\Y��R �H�M�~a-8��s�p����S��&���2Q�Fw�j3?}�x~�J�k	��6�V˾_S����ڠӓ�O#�H�� �,	����_��a�)
�sU_�fjgE��+;I��	g�"F~i��Ax���I?UbW��A�,u�[���J�Ir�c�)M��=�c���{?@�������Ƶ#�uJh�[��i눾�I����i���ˊ|I*��Y& 㥳E�V焗�~jċ��5����ڠ�D<�?-d���eK����N&����{lŢ����ۈ]*g�6�ϝO
 ������QDʘO�k�j����Lo�@�ǟY3��d
��1 B�hB��<���.JZ�?M�kZ$4� ���I�܎��M���m?�x<p\�a	S�bN)�L���Dr��Cs�Av��	$���4�G����Ӥ/]��_�~��������J��=��Km�&�XߤsZ����?+�[,�j�B�D�\~�/!�L~|ޘ+��q���1"G��c�k[Oj���;�N$��~���e�2aĦtm���c��&gmi4�_�ߏ[�&�Sõ�n@�͈�RǿOW����4�*
B������xNW{�"�KiB�V��*`��G�Ƿ��w�����TT�R|����7K�L8�=T��Y�`Z���(7fh�Y�� R6#��~1Z�X���.P�
s(D	`6 ����'���Lw	$�����i�&/F���������]6�V�ӥ��"6[�%ݏ8-��]�4|]��h��}�������*�S?���s�#��m�Z�}�!o16�!n<��g/�ޅX��k�.63���t�qq�kO�.�|,��$�lf��o�m�������UҞEA"R�;�<^�k�q<�}�{�J1�vB�ձ_��ƺ�n�O\d�5��j���qêw.v�2gt܀���3�39�Pg�Du ������,���U΢���3�80�/�!���\�gD =P�.�u��|�Q㘄���B������[�h���&F��`[0l'KH�Ȩ�Z?���q*�G��;�k�g`f�[N�)�I���-�,��u�?�p!ӻJV���T���2*��q�s'K��\=� �M���a������k���i�OU�x�SFS��^�']�hUu����2�P.�j0'����?K�"�^)c�펤 ��7���Ԋ��,�A�~;*{FN]�Fա��*���Z5uT�<�I5oMI1������_����w�0P �]r�0}5K	D����y	���*�*Lo߻�(7t�lD=^z=��8���;�R�D�~اU�4�A��V��4>��f�BE�_�'��yF¯Q�f��Л����O�_:ꔴKr������myvZ+6��!Jnf�:�]Aëc��s�@�8���Gh����&��RM�IO:�T��XO�%P���FIa��'����X{xڊR�K��{b��Z˩�mA{=:z��f�9�E��M�PNbu���w���J���F�S����;IB�B�B�K&'���X��p�[�m�^� �ݺNg< �a}zDb�!da�rd�3u�t
�E�����_�Z��ܱE�_NM0�¢�d+z ���p�1�ϑ@Y	۰�TOʨ�>�]�3{�������J���3y'+X�|!�9���f'�.u��_��R���S�������z*b��'յ3G"*��>�R�C����PS�!v �wXs�&4�
	���R�vvJ@�D�J��ېPGa��|eE�Oͱ�Q�ǉt�U�T6�3��l���aO�`��U�1�����q�a1 ߧ9s�4SYe� �V�z6���\���wn�F��D.W���0h�oyׄ~��������φ\����I)��YwPf
n�Rբ�:�5C��}�����7	�HV�\�<�t�7۶��r0qi8��'܆a����iU����^q���{R�qt�2s�I�3XAȺG��Cg��/�=��S���%җ�5�._?�fI�eT�V�{�l��)���:`1d�����"���7�p��zפ_�Y�̅������G��f]�O���������5���/w�Bu��J�#���_����P;vS��|
'���Y�z�T��9̞�~}��N��y�.	�&Rx��j*�C��Έ:��;�t�\R
f&yds�g�Z�NH�_��@�M3O�A�7�B~���C�;N�����#�s�>
Vh�|�t�ԕ?��6�_F�5��t��{��?iϣ����'+�qA�۷d8��D�ίG���5��b�k���G`�hGxK�鈫b:��YKW3j]�����qQIl�"V�6����K��w�=^H�b1���>g*5����WdX{V/1��2y������\�� �o���'�vzQ���6����kQI���;.g[�E��r�
ȥޡr4b�n�1�Hp!J��TS���YX�n�m��7q|;��+����}�z�Rʘ�����ZEM޾��ф<!~>�q��1H�����À���=�I;��	��ߢ�E���:�M��O������.�i�Z��d�Gk��������f��_�(��/�G���\K�Uq�B��9p�����8Mw	1��ؖޥ��Y?U&�N@��ۢ?z��eBGt�u%�|�=�����C�~����Q��/�]յ���w�����?Xc+0=Pa��L��faVkdU�+~	� �g�'�u�@!���#׫
�%���� �Oz����h��R}_�	�
��J�����vHsC�؝�x\�n���/���� q4�ZU�:�g��ס-��\���woV)�{��TN��B�O�@t���n�)R��o	����U��8m��!�����b�}�����/}�D�����Fwz��zL��VA�T����Yi6�P��D�����k1%��l�5�#Er�1<�R�;��j�r���5QZw�L2����Y�<��l�_��f��qz�� {f�6�"�x�ǫ���A�����Ԛ(\���Yu�O�Ji��8����}_�dv�@���K�m������ޓaz��_�ċ��!8w��b���[��2����ų%�J���
1ZS��Q�p�~
���Mz5�.i��9ZI��(���G�[��k�թU>�/7��:>��7+5���e��Rߚ����R���bN2�&Y�۳��#����ӿ/��[huô��в-�+�
ʒ=�<]�<O�Jﰱ=���������wiWw��
���Ԑ����$AjTy����`qB�wG�P�M��C9d��In,z�pZ�� F۹1�ߝ\��1�(�	j��E���9���ӗh%�n�z
=h��	��9�}��2dX/��8��X��{�^"Vkqfq.�
p܇�lVl�u@���R�Ũ���k&n��$P̵�����㬿P��u��s��[�hl�d����<���!�Rx�v?�)��>O8�n���=pI�k�	U8
J��yWH���}����C�^T�G=����fUa�|�����$c��m\:5
]7�c��1I����)IzIR5�M�#]�����2�2���oG!$�>F<����dل�"�Bɤ~�rx�4�{+��ڽ�
e	1�߹�ӵ��H����:{n��A�Y��OmP{�j�SA�ϴ(�˽�E��S��*�L)��q��V�5��.S��Ak�ho�,�Ak�`�j\���2z#e�J����-bٷ>�'v�*[4 b�_ک�H��g�%����ͺ_�+�)v�=�G��/�JR���
<�݃���>�<*{��0`�׃��K����b������)���y��#��`�U�9����~���v[�e�	��vs��Rd����������xM�{Q���֩f�q*��"8�5����E\��(8�����o}1�7�����^G.��3�]���,�2��;�{��3�/���݅JS"t���p编�@1*v"��ٳZr�`z�z��;�Ғ�޲�, #`�K�~��p!+�Q��b�E�����R �t��:H�A�ѥ�R�мe*��1�_�����q`ꪍ�e�
A��U��V���0"a����>�{#W5�p�z���-�@i4�U�����ۑ��^���;�U[�4���C��g ����p��.7���͐-OO�h��	����L�0'�m�Y�-�w��n��Y��2R�����
L�����	�[v�+��6Fy�8{e�>��:Tv�=fO��v�0��,!���
kU���}q�4��S7�Vh�#+u��'��e}t~4�@�x.��I��y�lt+U�|��a�]%��n�)ֱ���U�mA���;��#����lF��*��]����U𻉠؈��so3��i�� b�c�n��V���$�N�>��f}%�1E�����Q�L��Tg^�)��?�� �Ơ���e���t�</�Qqx�`�������>�6TC���S��������F�D;���Ha]s��^؀�5`�u��:�G��o�O��;�"���I�yXx6�<+���3) �'���:��y��R��^�:��|��<yߍ�d�1����(����q�q>o�$=YH&����7�vd�m��(��&6Ó�V��ƸW p��7Z�	}N��[8������泪�~��CK�kiֶ�Z�,�y���Yq}��3�oh���#�֖-@ͭ��v�D6x<R�0�q����n� y6[X�2ɼ�����$�[7�������P^������ñW����o]����qG���	)�@n��,��#���	��뚑T^ʐ���.X8'o��|f�?�5摄����%kibM�2�����R0�pP�<h��-�n����Z�]�1�"�R�R�l-���,|Ig�(�-���\�;U��l�g+�t��>��ٌ}�NEr�[���MY�I_���Rio��}k�]�DW�8]��d\�D���_ï���=[�e�&>���|�<��b̉Q~�'] � ��������NwC?3�M~�1�:���3�B�;�Eh��D� q<�PM�[�̍M��t�ԭ����Cm �y�J�:��_s ��s7b��v�H.L}�#,�A@Ϝ�]���l#�lhc>���?R5�vp�-iC�3@q��>���Xn�IX�bB1]�4���?k������ɝ���%>�u'���W;�� Q����	��X�].������$D_���L�w�� �ߧ�F�i����1�W�%���ʝ��?C4S�Y2��<~t�ˬpY�1Qْ�;�SjsU�3�#�T"����R( �H!H�h	ɂ~�V������Ӌ����u��fl�O�Vi|+Or
����5��p|x�a��b;��Y��T��
,��a�L�0|�H�3��o����B9�~��j�m�X}5؜��&(Hb_8J3�g�6���{sg�l����z�9����X6��L��bP�;:�3�:<��Z�}Vp���~q
\��71]�� :^g"�Z0s�i�0}!�Ο��O�U���=��-kR�:���c,���k�!��4[)����A�Ыl	U�LI,���°P��[�s`R���7{g�V�3��5�v�h�L���P�w��$kA��/+���A��]CxPb�kΔd=���)r��_��t���
G�4p�o����C�����)'���,�Ͷur(�5�:�'J���J�����`����f{QʣYS��K�?K�iX�c�Rb������tkz4�:C�c�"�!:�Mu�W��EBH��(X;���g ��Q���h��S��m(�4چ]�OM���15�J�x����s!k޵�=s>v'�t��:i"�P�7�m�f���mϻl��G��S0����eLr&֪���� O?��3�(�X�*~�x� j=��>�XQj^4��9��Fă.0~ �4.3�T�JA(�j����Eyv)�!}��m��OA�3i�;Pn����=?�i��o�YO��9����>��K�����OÎnF%���?����n��aàB���2$�FUb�3F��G�L�v�w�{���E/Q)k�|�P�lΓ~ �/�9t�Y�6�K�h@�E���� |z�Kٕ�����h��FR����^|+�I�f�~`mzB�ޱ�&��˄N�*��d�m1�bĕE�AOX<�Z����wK{����7�GCN�5;��	���փW��li��/$�6��Gg��Qx{��=X������q��{g�Rȏ�������߀��4IĬ�t��g{�p{��G�����-K���w���e,������K�ЌUWM��@v�/��\_ <���K��`N��BY�L�I?�ɻ� oT�}m�2����+I=
�?:tTpF�Ӎ�U�䌅�=�{ꎘ�}���3?%���(�\ |��f��i,b*�W�C�Z�)��̎CuW�X�e)5�0s�ef���ӌx[;|_�=<P/�E�)/Y-��u���e (ui�n	�D�*���R+F�Z��X�1�(�B���AƅUhF?�$���������/��n�^�Cpy�y[R���p��lzA��)#~ʉ�[v}
uٴ�#�lR��5��B���:g_ڤb�?�UNV��\'B�!�s�{i��n ��"�8UQ�n���T�A�����z�a$�2�یX{,R<�+ڟN�{AzC�c�A~�e҈�*�*}>������mI'k��ނ�)x�+�������($���
��1W���O�`���Y��>�24�e���y�~�`�g�����cfKT�����߻��P�2Q�Q�g^��� �<��RN���3k�Ǩ�NS����I�+ͻw
lp�^�^�H��,��W��Pٳ��B�I�tĮ}��i�JO}"��:�k�.|"�{�rzgE�aU�M�2y�oz����~�T���/��>J�,J�?�W���=���3g�O���O������6����<h����^;3�*���TH���R�7M铷��9�ڞ0�N,�J�0/��6�(`Zu7��j�ü�G�$2 ��*��E�aa��j�j��/6��>��1��8���>�	��N��QM�);�d5b]4�ĮIH�U�gw1"�Nl+�7��5��}��E����n�~I��^�}.�I�?i�P?��X��٧*H)��8��X��5WCM�=t���~�g}Goޅڵ���(�l���r����?ߥ%v�̄���{j�|#��J
49�`I��yld?e���<I�a*f�Ԅf���,UH���3�W�E�^[k5UXdl`0�X��ۼ��F@����)#�o���kk�ލP������(u&G$�l�@�_3�c�Aqn�L�[��L�y��ri�T�88Ì�d���"���O2�󗿀��߻���9eG ͙���!��P�Y��q�?YW%E(n�k��ݙ�,O�s[v����`�]��rɁ�x,6A>,DX�,&Ƚ�nP�@+Y�u_�ɣ�T	�~�S�\������	��o���?��$^5��'���k���:�7`Iv��AJE�"������C��%�+{���-<w�+���v��V�!����*�7�,�� ������N?y����6��W8���1��B�b^��$���Z5"���b�-�IYLǾiiʟZ�n"�����[mR�������n�O/ҝS�JH�^�Ke��C>��s^�Q%�	�2~��d��^{�F���GB��>���Y�^��h��*�;�@�e��2��ש��%�2��$�n�����MKQ��M��i��b#%������s���O�JN{�X���K��خ��C�tB�Z}�i&j*tZuA?����8!і�t�?�V9�ڏu�v�MMړ(L.�}z���ȍ����KG�-�]�8�s�CN�</kN:;F�0��� a A���\u<Z��Q��؂�al*1�o*�;|�*�]��t;������2���fs� P�%{��5:��}cBF�x劂ˉ`��`��Eڻ0U��	�VE�=��Շ--aA5��^�J7��"m�h��%���f���n�ovq�'�PM��J��^�1f�}��{*�|ٳ� $!�i���{�3�M�0��'�je�����'�,���>h�3C*ٕ��/��4h.�R8V��پ�]0{�JR$T�Kz�%,�Ր����>O�	�{e��aI.0q]LG�b��L#����C�bNT'����Y����9�k@�R��Uڵ"x����%�p1����)��/�y|�|@��ɥ�����Np�"��Q�g=�lڬ��%4�Lj���՗��� �7>T���;'�*��(=���PfO�eA��[����	1��ʢ�vR������B`�Jf2��Î}^���PO	I��3�u�u:�ߨC��4��ghM��E�xa�	!�LoK���'X ��<�'��1��\�N����\��v�/���oU6���~ׯ��BK�C+�$��_B%b7n&���9��(��X� lK���9�&�+����6�v6�ph�.�
�h�n/�R]D�|�8Y�'6�9��mr��D`��!�R�h���E6���O6I53�W�|_Iw����. Wp�I�sە����d��O�`Gw2v�����%�Pq`rO�8�*��M�����yGB")
��
߬�k��2$Jᴔj�
_�7z�Ӣ3ʍXS9\��N��qrz�3uϙ��l��&�j��S��GAn1�;����U��<�{��.�`�'���Z:��c�I+��I�}s���
랑nԖ� �d��v;*�+'�&�+v�V�P�|o��d�P��`@C]Ix���I>(�H��0CB�.4������o�P��G��^T��Ռ�}��\�F�a�|����Q��ߥ<��AZn��xES�!,Jk�E�DRc4�Q^�K݊f@��'�G:D�����mK��2Ά��/Q�k���T�Y�o��F�D�S��E}�����l���޴pUW|�4�}'��5�����7��)��CY�0��ZG�������k\ɛ<]F���Y�1P?>��G�������"6�������9HbJV�;k��`r�^��Ū	��2ع�^��dZ�76p��8�){ޢe�
��3�5P�k��/�2ԯ�bS�əǵ"��Q��'����`l�H�Z�0ѿi�0���g�|~����S��Q9��7պ���GK(�B9E�������V���Z�Q���94��d���%����A%��.	�ui��K?}�e��`���NH�E�H�\t!<Q@����d�,*L\��;���ni�"�&o�|jf.�ٟT���P��q��J�+�XL��ayz��Wp���*&���*�U�+��;��z��-ֺ���x!�+|N�����	(-�hxy�6�R:�b�F!�m�*@4�!e�uOCjWK ��ۆ��+916z�o���"&�-F`{v�$����p��8/2���Z��u2��Mw8]��jA�;|�5�����@��1�U�V���Ǧp��c
�̨�FŻ�v���u+�x2�IJt��`�Z8��0�H?����a�#֎hO����.0-��P'>���{v��U��o���MO��F�>��la�p]��(���_~��qC�;���e�'�m*d-+�+O��� ̚p.pmy#'E�(���F�w��%NA�Nޟ�M�ꡔU��qs�D��M���S�5ןy m��o�GFZ����r�4��Uc�&t��b�;��AM�(H��i-�{��j�!nA��H��* Ue��㾍;z�He�~��{�|���$)�=�~ �}�8���L����{J��f��J�7����F՛=D�Dj�z��/�2̚�'��f��d����Gu$��k��ͩ�Kr���]q9��{�e��da�s��I�Hr1V�f(�W�����H4�c�غ"�o����7~@�/�WrT��ieC]�F`�ȷ�4C��Cc�B���C�O�4e�
��w�g��]��aB�!#�'.�Dw��0djͻX,���f&c��8�}�W��f�F���u�K:|���~i#˟ǻV����Y8�`�b$$Dч�}K�*�����(���~4� g/K�����Ȟ���ü��Є�9�	O5-��#�j��BZf�y��7m��:������������E�:��w��|�Z]OAF�m�5�y�3$��Ґ��k*�Bʑ�iX} ��R�\�?iV{lI�4R�s���lWj��󥪀Ġ(�����֠3?�-3���?�"SZ1K���n��Bb}�T
��Β3V0�O�C��+���:�V�U����mW暡Z��dB�ʏᡌ�����s��D��6�ߺ��#aq ��_b��|�y�����A.�z
�UV������m��%K��v�x��?~����C����lȤ�Y� N���j�W����VV[V&p4�=��&��?���m�/�.����$��A���Kw����5��[�#��1�*J'��,�.�S�\��y���� 5�Yk1*��aA�z�d��Ы���c�ў�#���p6(��w�n��2�/ݿS�6Ȑa��: K�jO��{�"J���cO�����d��f����fH[�fb�`���]�U=�3f�n����J���妉-z�+�#b�X�Bk�Pt�D�#���Wm�1s�tF�~y>gRgИ��`��0�$��<o���0'I��P���~�0A�j�'�$ʷsnz���WP�Q^�AI�� 1f<�����J;b;~���jE��CiHii��@�poI4O�p��3h$~P��1"��틪l�皕��M

L�+��69��u�&�>$���܌����G�c�ڌ&���Y�=x��TI>���6o���Wo42v���#�N�,���G�M��c��� a�@�J-N,��15k5_"	w�D���ġ����Ր����J�Aٮ�s|w��%�.���A�KU���d[�.����P�R�:	��T�J�\�FC�1�S�y�_9J�#���;h�j96�0z}����E�JhwW]�'���d�sC.�NF.�~�=a�k�U�� �=�a1��:3�_��z�:�t�?!�&R|%v� �%t�s�&�˿�}32�d��ؿ���S��Ңi���ui����!�	����Sv�<&+x�(`nM�8�X"�G��4��JĀd�S���j��n�8���ܳ���
�-�ߣ�Y���� ��\|��������I`�#҅Y�qޅ�� M�����.jX�>��1�|���E)��b����2�b-g�̼p:�7\=)��w6����:Y�(}n@-��0��L!?{/<����LR-%��X�(�ˁ�^��+���q1��y�8v _l�ٮF����!�h�ݯiV�~Ŝ��m�&Pݤ�E##�4��I�%6�>��:��*���=�h0_
O�l�Tb%���>�)��%ޤ�� Ļ´ Q�jDHI���	t�,o�k^`�IZw�XI�"�W��+���h������:R�-P3�L^/�8P��}`�C�ؑ����ّ}���C�8����Be��W/r=�!���/���X�l!d=������P�H�[��:�jt-�Eݗ�-e
���$ ��kzta����>w�&&�Qm�|8Q�σ�?	�F��t?�'c�P��N�FjZ�O�3=��dqd�e���9�r:/��\�s�X�QY}⥔~³ʾ9Ks(̆�B!���(�7KpvJ� g�PB��i�\,�2#=���h�y�,F]z��J��L�R�f�?6g�ꋊ��Q@e��)���LU+�Q����
��Iv&���{aXw[�'��j�YW�j����v�mXt:C��B�p�K1�6��MJN����A�uP�W��F2�9e�^���Vj�s*NPL���H�Hf �X{�k�6�/�X+�Y�k�S�����}��������ly��V���z{[r��5��E��p��Z�a����f���/z�������ey�뎣.i�\��Z�9Y6����$D�����J3�9�5�2R�Δi�O�姤��ې�SOϟ�X�Z��A�jqV+����fݪQn3���\��Q��rk����B���䚟�����s��eϡ����^�E�G�?�.4�����?�� �`��5�;h������ �Db^25�Ac��oeQ��$R����癩D�����i R3%��m�ɄE�G������'�Dj�nk�Zq5/q|=H���M��k�F������K�Ʃf&�b�yXK\�ns'JT������t��6�����'v�,cR��L�=��U��ۊ�j���A����	Z����A8h���s�V�b��p<���9�Wr�a񏤉ڼ*8�`�����U�	oGQ���ky��a��з��k�� ��-C�{&[��(GǟKi~�hÏ��zL{F�,U���ܕa�ls�x�p�3r��f`�wɡtZ��&@�O y�Iћ��=��L$1o��{��s�AG����AN��|���U�Ag�!��$=c��r�[^4��Čs���KE����E�۽B�ک���A�t+���#rt�3�ػKj6s!��wUͩ,_BRid��=G�q���Xb��9��K���Cj����ە�
 w#�(���ՆaǾ��*�f���GN~��K5��T]
N@s�3�F��ƌ�piE�y%��v�E���EO��U��苒K6>4fhy������D&g����aղ�"5��.��㪊$CC3����E��x���<���1�=	<h�o�o%�$��-�$_�Ͳj4��ٟ0�ō�륵:�>�%a1"7֨�#�����?;q�ݬm[�Zn�0J#�G/i8vgj?R���{���]]�o�&�T�bU��/e�TZ5Y��CoJqT���JZ�G�z��1��<����
DKۡ3b�m[�]
zA�������~�71%+pC3����}�W)�?[�+����xt��%^�L/FAA���3�+���=e�Ut�.����UIRX�m������~�L_�6�D���)�o�<��ɲn2u���DK�^Ԉ��~"��#�k�K�~M��zy4Rt��ݮ]MJR�K	��+2�؟��H�  �;2����#g��׉�!%����}ϫVS����G����1��8N�ꥮa�9@r&���Ɯf��(�4K���>5��#~��	�8�]��0i\��"Nn�Є��'O� p�IaxE"9�ӑ�\V���������m��j�_ `}ȗp�tSE����T�a�J�4�x�@%��.�m��|�y��KR$��j����d>*�h��R�W�� �~�*�������*K�X��|"	1ᱍ|�ݯ�rTbZg~����<权�f,���1�s�t��,�)�}��+�3r;�nx��?�C�ldUV
]N�R��Hy�2u-<N�X��[f]\N�g������r��@�����J��*g��J.Q���5�#<��ofܐ4���Oe�d�C$������1I�L������Dd���zx��G�@�J���ۆ���� �B����S�,ZF�%L����\P./�~��2)n�z)F���T��S��C�n��=�k�<�� ��5����\����)�>����,_�z}|�l��pK���F6s�H«4��d'�u��=9��b��8�8A9�<V��ч^�r�!������܉�7��F����L�%��c��t�j�-J��������N>�����+�}���Z�_壙���IkinP��#��Xf�ն�+Y&�����Y}���g��Z��\k���)P�;Q�2h5?��Ց�e��
�<��s������D3��ԙ��c{kAվ*�Z���A�x|J�p��O��fV'�6�҇Sȏ(�+��oDlW�oh!�͆�a��W2"\����Љѓ���L"_h)�������Q���0��PhD���5��ӗ��Yy�v,Uc���2s�#�����`��ظ�0wQkj�
���bs�N�e<��S-:������"~.�'l{�>�	����` j����@�f}.�TK���
����I�{��oN�3"wW&���u��dAY�5�B��|?%6���g��?�ƠXpNK���Z�?V�W��Od=�H���|�a� ��ٹ�D��|��!vW䏴q��g
$Hs�C�O�492���K\s��N���0���d�?�1pK�Gm�ϧ���B��LC�؊�fr�%�D�w�f��w��F����{���M��$!me"���yz�F$a�J3�a#U�g0���l�*uu5�Nv��!�ߊ��f���*2:��a����%�G��;>>��������;X����hPcaωYn�l*zD| ����gݙa.��$�'�$��s��i��%&0�.{nKu�{ \kǆ�a	�֏���O6����p�`"�̧�m�����n�c�&��#%f!�zfŷ]�隷���8-��A�5B��X=�6����>��.Lꠅ`B�P �ҋE�b&��\1t��a�B�q��'ѓԀ�$���=A�5��ST�t\������ݶ���VcX��x��W�
r���2�4�?\�����L�kx��5�GG:9�� d,P����4��UL+�AJW�2�Ӊ��k�"�5��j%B#o���pTA���0�}l��;.��	�B�z�K��k��݈
 ��}���H����8�l�95�ʋ�9EJJ%Ҽ*<����P�u�R��˲�w!#���q���[>$bz���ΏS5�zUR�.�R{�*��$�+�@�b0"Ȳ�������v��U���Q���0I
�"i��/��bha�<vm%Ej:����P��poR���Di��t#ܼ��4�%Lˡ;ؕv����ޗ ��Tٷ����	��p�ũsW�K/���y'����X{#�7ا^��J8�����81 �Cִ1T������b"F�}���Ɏ�� 7�+}7�9fD	bD5sJ9z҄�X)·�ϑ��R�A ��c�.�-�)�:�m5�����䒂� cc�2�fS�dVR�i�U�G�1�,d�ÙL��9��e�	��9�V�[�{\I��N�s��h��������
U���g��K�a,4>�@h����u:���&��wsy�:F4��p���f)��A��+4M<�1`�@�1B@�6�Y�=x
�ܽ=�OF�,�Q����ղHWó�����w�/<�N	����m�uo��)5��:�l-\V����k>���vH6�b^����Z����=��Zg�:�b����=�I�^C�r�>��{�(R6���G�7��Eg���8��y/�����"�y�ns�+�o�q�L�ʿ��+Ps�D�@��L����t�,�(��Qᨻ5ߜ�o-N�eW�<��������@`�y&�f�/�b��u.&˖�����L�bA��1\ �h?hO>�h4ǝ����N�H0i��Tz��tz�CuD��l�A2ط�b��5;���y�MTߝ� ���y܎q�7.w�L.�{�$�3ģ��jږ���+��ѫ��Z�|�I,���t�ђ����'D-Ac|���`�$�i�,��\Ҹ���Q���yW❴��E�X�-@�\�Q���1+]�P���.Tˆ��0�>˪�\����j��:��`�#)k=[&���p�kD|�3|�E	��V�E���a��]���
Y)y�V@�U��c;S/җ�Щw={�����8� 5y{(�CX�.�aZ.P��a��ʏ7�������)��T��W����2��+?]���^�F7ˁ�lE6����m�x�EyV��������-�Գ���o�&����������$��� X�1Hs٣���C�|�yc�Q\��`�.Ĭi����Z.W��Fo�1C܎��k�ȑ�<��A�Sꯁu���l�������,�ܚl��^�ߨލ���8�x=Mm����p�jِ�p$�\\�ل��D��cy��;�=�|�4(q��Ĉ�4�r��-mw��P�b�|Z*mC�/��iu���96��o��U^�ײH����x�8�n�y�OE���gꚃ0v�\��)6&t�E���;�x�A�)�%�`;�L�E�6�U3g�2R}�^��`�ʭ� y���}�^$�c��]�B�����S����8������f��?E��5���V���=H���<�B�k}�y�H>nŐ���d;W�F�d�^P�����k7�D�,�^_��ƕr��O8~��47O<g�\�W����l�ۼ����Dq��}\��=���	�ʰ��ܸz���e�8͓��SL�bQ�Z�iҥңs�%]Xq�U R��Uי	?���/�w��U��V����OG6�+֚0��G5O�o�j8�R
"�!�L����EoP��R[�#��(���>�	^�Ý=�ͨ��j#�pm�j�A[�"oV�z��vɚD�s�d���4�l6�$c3����In-�����������6���ۑ�h��M� IinF�B��\�ut�:�zҡYyz\�Q}�ޑ��y��X��d7���� �������_��/��1� l�5�>� �>fS������-�6�/Y�_�p�1��%фW�i�-*�r�ǥ���V��O��0� nC����������1]r��!��6{����o����t'�L����8`�n��ʆ�T�W�|��]�2 Ĳ�^�8s��sHXny�h�w'���9�C[��c"��\ �ӭ����� �j|>0 �&����C=�hW%�6}�*1�~��p�MF|Ɨ���↓SFt��2��?[�[C����D<114^��X��G�~RűN���\ߎjs�3���TD�h��
|�.��U.&� '5_ͫW�$V�NK��g[���L�r:��ݒ�Yh�tC�A�IweA����&�|;�c���I��w��q*?|˟3�ǚ28{ڵ�tC���P��5W�ʂ��H���\��8l�S��]��c��4n�/\:�,]`�^�E��R�u��$�Lr�Rf���|�hc�ԞF�R�86)�['.��	�A��0�(�G�_��v�}v�^��2����(����V8<������x�~����l���>�$ڡ|i����귤\~�&/��A)mDޞ�͏u`��_�"���ȳX&�1󸜷��[�oAD��m0����YĔY���nf*�.EID��'���^����N���^>���3^_������D��z1�u窈m���� �BN��v�k�ϬZ��E�i��2�w��rr-�a8|y�S�W�ab����
fr���s��X""�/���wg2�g-��X��iY�^bR�;�M�j�u�c�햴���ȑ6u�@�P��4#��'ix��?R!!;{B�U���hn��C#�[��M?m��K���>�ծE�B�ߘ�9zh�_�P���Ȁ��%J��A�̔�K�T�6rfOx@hS�˰�.�Fy�t�zB���3�&^����t�тş�Ib+s4��E� �Ä�ӯ��̅~��ʢ���>9G�w���h���~�zD�C솬[��`�ܛ�_�ԥ���<��
V��?E� �k���Y[��>U௬`���>?x(p�8V0�Y� ~��*N�<N�.��gf���r��yA�X��-��Z��>`��џ�fQ&Y��X��_r��0�.�'6 ���Ъ �2��W�6�f71�毭d��,y��m�W�Vlr�̅1�$�}�5�ݕ�]%��8��2����V�7�k�1َ DBr{����9� �/�?��	ݝf���z�8A�d���aV{��qW������a�z��҆w���rd���t�~���2To&��f�5�q���-2T!ۼ��[��U��e@�
\��/�� Wio�����P���K�-�74��o�vj#9�<kК��ث�x7�9�&�'�����Z3���R�P#(h���'��~��U��!���n9�:��7'"8E�I����ǽ^�H�'�m;�gy�-��j�@F���A����#u���SM�,�'�.��,9����I����τ��Bi�l�E��K#�Fe�������m�� u��0ڌ����#��j�Ң���{����9�)�.����&7�C�i�@�"�����2�k��HiͪG�-�˼s+/p#n�15�b�Ɗ�LD�*ǒz��>�ZI+o��U�`���ri(�-�ݿ@ǧ�?����6�Y�g�r,.����֎��$��m��qnw��D�%ڈ�pK8v�A�V�Ȭ��;r��A����+G�hr�kh��R#v,cI�/�!�H����L��I�&?f�Z>�I͈�!��/�%��������#�Q�bi���	��`��N��N��^p��hXM�&�~G��(�j 0��֣v8yqA��!�I�=9T��/�ǭ���h�����q�=���bڼ��j���WZY�zq(���h<��~[���%��]F�Bڠ53����-a_�<����dnݺ6�kb�G+�~�2�3��*4JG�)ߵf��"Z=�����F��!;T���u��P��ӝ��]LZ�>�E�T���vPT��G�=�
�]}Uʙs�kMh������$�l %O
k~z�$1�!����i�zk8	�RK"����~������A����EF�3R}����8�0l?O���Q@��H=�[��v����)n�(�=�օ�#�F�h�ְU�(�F � ���(@=ι�O1�h���$�N����q'G��*���<�����3�����H�-j��y�k�H	S������u�,ip�o�o�T�@��;P��AH�aɶ1���O�y~Kd�5(V��R�`�x���Pc��i�w�~���fQ=��{n�n����N��Ma�[���9[������x6,L��:� �R�*Gg������~Y�ekZM��a���%5�w�o��/hU1�".���IBڈ\�(G��̇o�l֘kjd���t�C4�uoF�F���-W|��bWlk1�!��a�����Y�#%�G��e��)1{�a����~MK�L��/�Ű�rh�I�TU��E��V^�lq�b���]�uje��S�e{����Em�[��7['�>]W?���z$���;�X���3��M1GN��]��+t��gǵ����k�:\�e$L����oTG����15������n3�	��D�Չޘ8��i�hoS�a�bt����g�[f���-8�@ֵ��S��HG%���$T�v?����KX�F��Md��O�WG��hg��`�aaCY��h����Wg�0��_�_��s�_;k'��=����ĞF%ԞY��:��)��ĺ.�<�d[ sr9�Ɨ��*�x�`竦y,C\c��B��<��ʹ`+�HE�Ъ�ng���'X.(�`mLI��X��8y��F����l���RO�٦��eV����8]#�Z�z��G�ZaN�}��
W'�x��T�	��4�ۖ���p��[wZnE�?��������2`5@9�Hq���J�:w��pG��Hف%�۬�������D9C%��Α����"�^�����)y���.�c���D:��x���փ��7)$�(-����g..���s"N�h��"b[m�"����v�g�N�D�f8�L�M��
�R��������)Ј���[���c���_*��y�e�in�����l*}z3_Z���=�#46%K�^�S�
����B̴Y��7��Z��o�wf��t7r��K�֖NA������=��UweS��a>��n���Y䄁!d	�My���&B�q�X�>��xQ�5���Z<�MM;x5_A�;cq��ww �D�N�m2�p���wa�*ݙnq��"��[
�w�a�XǠ>R(L�C��~8Bk��P��C���l(�=��I�'(�S�^^JA$c�"�W�c��d�x	X�A�:ՐH�CHPa���%���k�J��Я�G|��)i�sW�=�/������:�	�����:�%D������`����y��T�
cuK__�:8~qC=x%[����@e�ȅ�5M�f]�O�ױ����A�I���jP��ȔU�b����GQ��mr��Ы��0���S�MY8���a����@k�A�t,t��'O�/��Cbi{Xy�P�DadG;JKT���{��ܨ��3-a�x���+Mb�dI�UR�<����2�ur��b5��%�׆�t���c�+3��Ǳ�?��x�1�A�1�!���?�D/5���\�� m/��ւ��7���\g:?:�+��lc>'kȉ��ȴ���|�ֶ]�`�	�N� ]�_U]vq��#}�׋5N\��I��><0�q(��N
f�c�^�C]rH��d��p�[�Uj���;��)��㸑��f	��ŝV/W���O}�*b��Ze݌��$dE�t]��`�q���&! ʻ�MO�׏�(����@=�n�9]�p�:�?�`@��v��C|���ʥUc�$��s%S����\��xa1��9���O	w���uj�����"8;{����ƻsώ�{P��������
�dS� �x���w��tM	�����z	����N��s��G�a�����偄���,d���g��b��z#��f�X��=~!��������i*�P�A���Amd��.(��4����� ��䴼X�˧h���(<@۟���UW8�s(d�8�8"�R)v��@��Iʣ|zlbV����rh�r;�S���ꨇ:ȨHdr�b�%��3� Z�'/}�&�/i,i|]�(���0rf�@A�����3���B�A[��f�5БU3���]�P���d�#�n������Wd�;�Q���I��z�Ζg�@�A�f�F�?��AmŤ��h���ܑ�4�bR;x/�	�u��DI�v�؛n1��8�X�Vd�S���x��r��鶅}q�pv{�K�����g�/���B�wi�s���z�&�� ����l�(2��̲>�����JT�p�k	���{�Rܺ�z t�(!t}�L]$�6N}��=�_�W���V�B���]�̎���c�ڣ}`���Q��h���HQQ�8L��t_�P$�+i%Xo߀w^��t){�A��
MO������Ͼ�A,�LQ{@�AH��8������U/o=�-
S ��D�q����3w���[�`M+8�q���Xv�� `Y�`!,/�T��[ ���:�������b'Q�-�+�Þ0�D�{&�j�d3ݦ�\�h���o�|<O>�YU�+����<��L���L��ҳ��8u���s�����,�!�㘾�]�ce�0�%(�as�t�wDh��q*���s�9��!�<u=��)O��U��TF�6j�b�
>��$/�!W�Q�(���轅@2MK��N��zv���D{4��ga�F$J�u\�v��,���2][��D2&���]#�fѤ��=�J͇nT�&���P�#�ʃg\P4E A�A�9G�F��3�Zq$h��a�t5 Y�
�)�[��׵��V�,��� ����=�o3���$��
Ry����Q�xU�����Zk�UѲ�2�.�����xc�j�� �[�r�e�B�Tu��{���,�傟��/���+���yŦ���ik�&Jmp��̖h� p��ˠ�mX���a\� j:(�)	�c	�d��*..7��
58q�Kzn<���yʫ-�F%�8*�����	2�4g�	
�_��:�^�w����;;����:�87��t����}�w����I�Oxw$6�D`�v��h� �%���{A�:���D7gM�s�s�ܝ�9`E���>Ͳ��.���OgxN�[l���t==���E��>�!�>!���f���� �P�2r˂��ګr��5��BF��~޵�8�b!�0��q*��8�8��i�߽�tgE�Q�ȣx���v�ƌ���D����������_���jBn:�Z-�n��A�Z�'�)C�.wjM Ȟ�<��^
׹ T��s���>󁧉�#��-�����HI� `>0-�S�2���彫O��3S�I�����pW�b��Dt!b�*�8�^��>��+�����[k���FDo�+����Z5$X��U@�u��ϛ�/U4�Bq��N"Ԇ�+����r�j�O�^Eh�O�%�T���u����#-✼,ʜ�s�S���N�2u���hr";�8_oY����Ot�i���M�/�业�3[ �?��#�;�S.#:�ȭm7�=���s`��_�CY��s��	���2��1���o\SS��J����_���s�����Ce�_l�b��qTl�uAb�M=7�h���R�����~���!iݲ�7�_^h� �UYʈy��p���C���O�|�$P��i��r��؛?�*
4�*�BuZ�8恃ҧ�u�) ��j��a�9sO�&��7�O{��$/��QT�3����8�p�8λϜ��.�N�����7yy4�o��B1�6|0��}����0]KN7)��4��f�ŦT�eh~^�E�p7q�'��OiL(��\6�O�K���]����Y�1dc|������p���0�a�GCHKB�f��Ц+�T1:nqA�z��y�um$EgݩE�>f5�&��;���GS�Cޞk�H��~�%�����y�s�M	#/#P�\I���eo� ˑ��D!�U����f��|ű��������A4�teɟ�eAY���[�n�����k�/�2h'[�>�-�k��s��̗��~m����� �a9�A�pkD%jR�R-�5��W�Z��܁oF�<1���lPa�a6$��X~�����y�~\��A#W�����Y]�(]K�-̱�zO
�����sz`��4<"����^��5���[�#�T�PFNZB�,CL�so ���r��td+<G�S��b���?�,4ޟ���N����� L�E=��X`��QN.��'ۻ䁋x�	?	j���@�Y��x��X�k��Ѿ3��[I�D��#�3��*��%��E��VfJ�T�%�!��twa.�1��X�}=�'�QM�u�Tv�#n��������%1Ӹ��t]�\�Q�B�_�-�(g����v0�%��(ҥV�#Q��Q����r���z�Q6V�~���K�%�2����ҟ砛#f��y,:��T�uV����vy�V�W�J����V�IQ�;�"U��q�]6�~�R�J8��ӧ(q�W�l��
��K�%8 x������ղ,M�&~�$<��Au�#�&Ύِ�M���1�g=�|E�S��.��lP�S�W/�"��B�[�P_h��U9t�7��L��.�0�o��.(�+\ ��p�t��S���g��*X�!��>�w�èX�$�c������Z�����^E��q_�.��KN�:y(����I��A&�y�9pCk�/6������J�f��:m����F�^�a��E�Ar	lJ��S ltx�����cGک�&�����p��"}��*2�KM�^�i� S�~F͡O�GS#���`u���mm�'&���u���D�r��ЛwN(��te�� ��ӄs�dm���ف���cZ��a�)nV��f���@�ɿL�Bq"m"��Qڇ�$��rT=g?��=�����%��hK�WU���JÊN<$�5�x]%N��>�[��4��P���_:ڌ̛�����i�;�}��3��w���!~l������!|srt���������$��qt$�r&l���^���h�*P���<ώ6�6ӝx5��&'6_��S�Nc�= ��6�Ms�2AY�)��`��}���7���)���pM�U7��y��k� �����֜ש�V���r0�K�A4�Z:ݾ�^HXVD��8���2Q�
	��a�ծ�p�����O{�t=CB����Pmx�o��!��"Ѵ����@Q[ӎ \.NNL#�x�M
kl1@���L�W�ү���0,sL8b/=��Z���b)�$�@#�C�r��H|�>��t܆ Es�_i<��\@��UPX�ׂ�.��ݙc�k*
���Y��{dJ���F�=�R�$�yA߫� F4@�g�C�v�(QS >��w�)|�xy�{���Ҥ����]6%S߶e� �r{8��<���:O�zlKX�-���Z��;����%;�h�k��H*���\��p��<�i�$��3���暳R�wToP�5�f+g�O'I�)�U7�)��C���q��y\d�3�c�Ռ�1dfH�;W���[׋���W���6��;a��d}�N�� ry@�y�vk�=����b��'4���L.$��Z��������h�<��=&kԕ��e/F0)CڔRm��黎n5
�28B�گį�Am���5�>>)�@�P��#q\N�5.�,؟�k=����D�0wCA$�߆]w���
|t_�|��-�CV���1YUp��晡�oćV��xc�<�"G�(3vF�d�D��m���]�>v�>�{|v*���;◒�-)��}�Y����YKb댼�)�{I�Ǥ�N���Z�.,I�s�avT�TM�����m�GPΒm�Ǻs���T\4�АE}�KVg ���m�߯���s��6���rg�%��Z8��pǣ����ڠ"`�3aV����Bj�ptV'5��fE0�Z��7�����æZ9� ������ ���Y�~ǑǮ��ƍ�j�IR��G����{d��7�̦�;�
����(��nq[�}�En\�¬�?dO4���ȹ��f8�b�:ԗ$YTq	��	+�>]S�����l��/@�����$N��ɳ���"~ZҘvC�m1hR�u�TZ����E�N�{c���R �Q��S}�c��[�X�+)mp��t�'r|�H�}v[�1h*�~_�s��8A䝏N6�l�Q�ǔ��>��*�֤��t�D6����@��b)��{ރx� Z#��ǘ{�e]���P�G���c�%̖~**�{�sB�ha:�	����Ȟz�:�e��L��;|VR�^��D*�[���ɽWI+vc��c��z�N�i���'�*sJآ�3S2+����ce�^\̀���ƴ��,�t�N��ڳ[簹��/�����l��ewt��E��F�]4G�d:�%U�Gӎ��-k�e�t1毪4^&��YO�- 
�::?f�P<q��
��#g~�E��y�)�r�w�9�>���m} �Y�zF������Ԭ;P98L,/NS�K;mI�mot��,��d�63�E��>�w��a�JB0��z���f&E�#�8�Ɖ4�lφ*n5�h�a���Y��݃�� C)&I�&p6
ˆ���<���0�(Ӱ(���ނ��	���i�]��� M��C��A��:����$��dK�:=id[�5r�x&9(��p�bi2^CA��S*��&�ѐ�1	��Ĳ3��ZJ,W4�X�_�R��v�+u@�p6��M�6w]�F�rŇ	r:�*R�����m�7c�+�d>]���6���2͹�p0�Ezf��m��3!���g�v�DF�_��z�L1����P����=8��i�~�*gM�����֡�8�}s{�v�\�.š�\��Cx�1,�v�d��̅�*A��0*��6o���&�S�ؖ�MZEΕ:�"|ȷK٫'`*� ��b)P'���A/b��z�0vgSt,u�������uK-p�pF���z��]���O�7�����yб5I��I�֖����r��,��Մ��/mU�����Ћ��U��Ǌ9'e�V�a�#<�s�31�2ݐ���� ����	[�����꫕���=����0<��(9��)V�\�Q�L��$��T��7:d��%�]�B(�&iٽ��:�v��a�<	h�󺄛��Q�JV����<�L͒}8��ݖ�:�x����ڤfrb{>�Z���}�>�@_��9�����4v@���tN>��pr��)ެaa3ͥ�ӑ���ԍ�\b<�a��(g�C�-&�,Dja/E���iP3U�'�P�|���Ўf�%FI�/ѵ���HS� }c��ɡ���l�0ەɟ�(�;��B�F@u*�O��X��D���`I��49?\�	n��N�0%��Rq4~y�C�n�Ls���`�	�*m�腰�Z�������P�zh���e��dB/:T�i�[q�7V������z������@���K�xXԔ?P�zY�[�5�ϗ�.��=Z�7U�Ry乿E��|k��W3�*�h\Ly
qN;S-1�X�S��_y���q�-P���,*�"6��8���5_�kY�@�����r���[=^d�/��&���𓹓�h���~�����gS��|D��Ok�Mb�����)J��a�����jnE��PC�V�MK
�U�y:�=a�B3�a8�#7G@�2NbǍ�J�8�pt��{3���C�I��RYf<��P�d7��%UM<;�^����l����a����o������|��e������{�����&��c�k��j����'��S&/�]���#*�Aƍ򱞗�SLJ�8ie�����	�ƺR�yg��M�cL8u�V�@�#�o�I܁\๨�B���j���.)ՠs�WF�]��J�:ז�Z��ZC@2�;+��C(�gy���\��Bqn��sq�<��^/5vU�;�ѝ�!\��Jf���X��V�"v����Q�Z��m���$ME���\_�.��Vf����8Fz��1n� �z[����_7-P�zk����#ﰳ��i1���|�	ψ���D�$��6�+�` @G��8�?%a8{�֦Z�FRl? ZP \�-����y<�N�3�Cb��I�7��1<�� ?�oC��6�5��#�g�y$3��[��w��TR���T�YA]
������Ц-^�6��"��O����N�n���:Cy������ے��IW
� �<�U7�P ������	�kQx�`ik�"g@���S�U�2���|}���i]���}-�N�����c�u�	�o���Է9mq�W�'oՠ��Zr��L��k�񞋷a$v�4���,��d���t�������q��6���I}�:�߉�}�XQ}}��hL\��#I�ھ������0���2���*8�h��$Iym�?X	Y:�]��7��5=�PP�T�P�le���M�����[W���A6Á�2��r��>�nǎ�k�	Ǒ�I�������/P�V8���@w>���,%-�Y�Y0r�ʆBh�%�N�Sq|�^��nt-�?�!ˆQ�Ja!R� ?���������}��7���;l��B�IhQ��{12�p<����}�.�9�LQhgZ�7)���}�x ��#�7!Q�fRo0<4n�N��
n#��Q��Aa���(o%P�v~|}�yv�.���3U�^��L��Kx�n��9Q�ݎ��8�9y����C�7#�NBV���%@H!)���,̫|���b��kp���i�M�yR�`����鲝Vz��Y�W�x?l�=Up�4��N�XY.����Yp3��`��gW����=ꘑ��}������ᵬ���J��d���5TDd�M4B=���QT�cc��^�+�	��1�M�%�t��x��$���آ_nq�|T�&!�OC!_eH^<.���\��>!Yp� �}#�g��y)Q����v}T��]�n+;���6�k�A�i{���l~�:���5sc0W�]�N-@�ל�m�ڥW)*� �BF����իy/������ %�4����Z)�����߻v)�6�z��P�mF�)i\�V�/yQ�i@��#�@q�~A-�ߔ���a��`\.�g(���(�s�4�O6��g_�k�(NN;8�����1�������}ń��PR��K�.hYۚ�$�%�ߧ��q֧��O��A����)(�Ua�J��Ϧ(�z�7ni� N{t�[3�ٖL�3'$��dO�θ��	gq:QrO缤�	�׮^�1����+}E�E��5xV�pK�����JiĶ��� �L��!l+�!M]���Apn���^*ƬN
Fc�����v��n��.�8�7a�pXM���v��*��\]�'#|<�'�Q#�VO4l�� ��]u��N%d��OV�Dz���c_�|�R��f�;����r.��M�����(d�����*� 	:���̜��ꮚ�v�N��Я�d"�g"����5&��;��c��<��ğ�5@go��qi�K*F}Ç�WA�lٴ`�y	L��p�[���M��#�L���;�C�B|�6�����4w<���n4r���	��3ߥ�W$�x�}_T������	ϩrj��^~l�V���5?&
ݼ"Y/�T����CF�EP쭏
�n$.�}�[M�6$E����{�����v�զ�Ss
�w�U��ںo�br����/��"}�u:�c�:���|G^�(-����I��E@85����Տh� �E�5�O�rne���ti{׸�)l�X1� /��Yȳl-�F[*���_�+�pA�'(��'�M�YG���4k�T
F�543-dUt���F�XK`��>L�Зz��d���@:>\Ʀ���Ӎ����JNS$�ߺ][��Y~���ֻ��nH�L���h\��� I�Z؉�^�CS�.l�i
�W�Uth�<�t���o���k+
�bS�<.�@QE���~
4#j�I@�J҈qr8��ʦ��d�g	�.��%dt�A�|�R������zШ�j�����v�s _n�Z��m���1���=�0Kܖ�z>{^%����ZB`��>�5\=�����`ke��-2�&����,DW�m�:�ldbC�J�[Y�̈$������6��:��(g�k�Aq���QIK�aWK�#K�K �h��1����z�H *RC�s�դ�~K�xQ�	�P����p��q��'�H���ak�;j[r7RTA1N���F��dV�I�{�!ڋ��?��Ծ�}8*�3;6Ù�d��+�����+o�k���z�H%y�7��x�=f!o����W��[e�Rߜ $��d��)B	����@�\sCF#�-	��T|�WkNS�%�P��y����ݠd�#�ޏ]�_1'��B�ޑn�%0;wUAPn�(�!G-�] �mГ��LwB�>�!��d���BW�?�Ѝ��aX��\��S�,^gE<�&E�`��@�t~���r�	�M0V� C�Fw�s%ٓ����a��2sK7X�r�����,����rt�h#��h&X�z�:�.0lb��לͿ���V����W��E�E�@ʍ�l�X0�&��#�sm�M�r£wU���`�Y�/���j0=�����@�����A��+�\���t��ھt�]>�0�Z���_"5�8��{��[���Sç��W�լ����B0D�r��dD�տ��ϵ)�D̵:���X�g�^��������wK.n�J�[�հ-���18�F�P�h��Ȉ�;<�^���P3��Ml�����m:�O:�O�,8��@	�ij�78᫃��$V+`=1ѓ�[��Z'v�-dXS�����o�t������G����&4��+�5J��� �'I�S5ߞ �{~�j�0K
'^[�N�zk�"��>	���%|�!
��%Oa���0r��OƏC�!r����
,��F��<i���|�Qu�*08���co���j���Ɖ�; �/�az�Y-��ۄ�5�u!����$�N=PJ�q}6cb��x��lP��U�L�N"�,�:�tJG�E�!B�r��v8D���k�7[�Z� r���I�KKE}*�$��p�_1�}|�Zy�5����b-���F���i��۞�������{+�O"�j@N����`���^,p�SS�ڲ�A�&�C�s9�xb3�,��P=ΏAپ�e�ʅ��TR�8gy���4yOii�_�-��߸�ހ��B�G)�޾�$�3�s ZN#a���� �($�NX�i�x�5W�B���9��LES�o��V��<QB�V���j3ej��'C��`�s�Z3貟��7���yO3h�5!iSc9�����G�O�.�����p� ��t��a�1�4���R<�@U���&"�c���w$��mz�*���:�����Z��Ղ�Z�}
.� ���t������ւ2�xn:5]�^1�V��"�cp'�{%顗��<����i4����	@��n�*['?�=:��5�y7�;��nxP�ey��5S�~��|� �/Z_�1e�Z�C/ ݣ�R�~y���F�A, �H��i����:ҋ�a���2�����������r�ڭɣ��/�2�Ƣ�ܯ��/
��=��'�	'X�c��䓽7�=��O��$E���=��jЇ{��IyLu*�pW������L.ȖYt����3\���BF��%D��qZ���g�o��~�*��F�j_tN3:�Аozf�ou�c-�W>@bT����u�x_S�h���lE�+����5�OШw7��ˀC�W[���ř��~A�6D�t�g6�n�rɐ^)K�ћ>�a1L����F���x�Ҵ����� MOSq*�4�+8n��mf;cR��4�c;F��u�3����E(�:��A@c�#�3�B\�d	�#�������f�v�BW#e���\�'�c�)�h%���a�D�^�+�J)*��↫<�'��E歹XM����	(���FMs[��
6��� -��c�Qg/O�m"^=jmF8�ژ`�8�l_l��.��:^R��Ӡ}RiQ+��%��q�+
%���Ǹ��P>4ȧ_k]Su��u��L2x(��p%xX�j:�� *lLL��p}.5���C��p�L�_��X⒥�J�T��ez�Z�l�rK���wf�����v����OR��y��ބ�X�h�1؛ �ȓi쩊}���}�]��l��zb�<���euЏ����D�!���y����]u=�쿇�eͳ@��C��+E>�hPa7f��s�{ڹ����g�+f��1@�B?�X�}ϗ�*��t�t�w�S�,�Tg~:˾O�������Lm�X�a��w�h,<���Fo(�4����@g��A���h(��g�_��R�2�������EY/���	��h���5�+��$�oӄI�!i�����#�v�Yb&�+�G�(pL�^�߳e�G��Z%�Y޷��^�a�z<HHi���b'I�-T���4��{��C�Og3�D2Yrg؈O�s���j�*�I��Xr�f��)}�f�>��C�#���lx��#Z�q��]:q¦.���J�(��]��o�{Gx�S���j?����lT'��0U�X��0%�5���#������'�������/�}�7&T��D�09����uY-ҡՅ�2���X/IÍq�[�
��&Fj��I0��l��λ5���!��kz@�<�%ƀ��ߕF<��%R���T�r:��0�t����%$�yf���x��,oU34md�����l�r��	��o ����2��	D�ܵf�V�I�Վ��5���A�W��n�i�,l*�᭙'~��,�.��F@�fQ��FC|�z��T�m���$|`�t�2��o�ѳ�.z���ǚ2x�N��M��B��S�	���a�G������R� 9��1�Fe�������I�c�o3���+��߱���j�H3�ZցQ�z���a��(4��K-V�89�g�N���}[6MW��e�D�{�#���`w��а�؞!�Fo����PJ��r��`��a�&Y�75���Fڄoaf�g6�C �a�nvkg<{��*:���A�ϙĹZ)�o��?[���Z�,)��˾0���홇}c�ZT�3��]�15<OTa&�!�.�U�0�p�?H��{bB��CtFo}�jۜ(5�o{?~���o����N�gPL3�pw�*��2����ҳ�]S��w�C��F)��hk���C�V3τ�I��(b���}0=�����^�ັ�r�����	^��(;��֪��4�K��-�:��f_� '�Wy��nc�D��:�@!	o\:n��]ΐ���Y�J|�Ǳ�2�l�5��������ɇ�RW�_�f�&�>��kJ{���oWA��$���N�bT��.�*�H����l0����0T?��5����8�W�7_�ܩ7�1|G��_9W����ɷ��3=Lr
@3�f����}s�vкTH"��?�r<H��3�E��񀵳�s���;q���O��m��EA�z6쒅��P�$D�?����z��S�s���X�9{DR l�70���+��������9�:��X<��6��@�S;"I�y={t�@kYa �{��$�7i���Z�΍��P2$�Z�+<-��U��Lb]X�j0C�	*3���l?�S�#T8��`�2t*�����Lp�9�G@�z����X�r�����k�^UV�u��p���2T��v/���g��sz��V*h����#-����e��=.�k}1� �:��7�ס�Gxm~������QzX�W��?�b���u^����vǫ��
~(!�D�m��M���e�N����՜h��� �/Ư:�*`�"��"D����l��6�e�23��<�*և	GAϭ�g2F�^�zvw:�g>��`1�J��[�m�e����Bɡ�����X���PjoA�5���-�(�;L}5@��sÛo��@����߾����A�ً��x拆��B�~G���;U�,N2���"��i蚃�f���?B�0�썉+�"�����f���CR
�Y�εhÀ��һ�+M�K7�#ˆi�kU'��q_@9�U���I�=����+��{���gZ�9�h=<��q�;���'⏠0{��kѩ����xt#�M{�C1<���8�ߩ{r�����$�� �X�<��3\���b���,3�r�=�|bh�V�_\��_���b�T��R�#��3���6�5-5��
�y��0CM=6�ܛE[�[[�I��B3�1�ޮޅC)�����>@��=��� 6˚@�4�o6���v�����!�Rt_-z�W��\>��� ���!`�n���)�j�V�I��B 5mo=��H�������GW�԰M�߯	*�Q~��y \�e�m��g������*�us�sk�R���K����'Q�F�0��͜��z�E)lS<�t�����&��&�G�A���>����Jv
�?vn��i�L�=���[=s���>'n_;�잫9�1���+5�O�����@Z,M
�8��k`�%#���H�[F�mnȫa<�1*砇ƾɻu�a�����ugI<u�����P�uo�r|��Ri5����|x�����W�|��&Κ�_A1����aO`k��m�"�O@L�k7Z\�*��<�W*���~��f+�Pe�(��Ld#^�y�{�ң�������?�\�S�8 p�>�1��}MK1k�}��d�2�pXQoՍ�6���KU���xǛ�����31�c�ۅ��
����6{�;
�7d�vz@
=�Oϧ�#��hJ�W�[ �X)ɥ,	� ��s�!�ʼ�'��xȓ_�׶�D�V���{M��ϛ`�e�,ϔߞY��!*�¢��0sܓwg���+7���A5��T����dS��uJ��sL]$�C��Gs�|�}4W���x��w��H	�y�V �����f���!�N�J���)<�C�.�,Iy�>�Ҭ(�O2���7��"J^em�p$�@+>��86P���7P}�<ň�%��_�b�$���6�R�/��xW�Z�\�/c��	�uG��?��e������'�|��Yb�搹J�Q��tt��O���,�kW(C]8�R2���(��ӝ@��N�E������ͱ��&���cFR�����L�a��{PO��O�.XG�i6ʁq2F�k��I��PR�on��Ԕ B��:!B�#������-s�N"n���Q��.�٤��n��J�2^�!j�%�������Δ�žXAR�5.S|n-2^U��RN71#�
�w��|���A$���7���0����G���}�"PFY����t�+�1.�B-ڐ�i�fS�C��rN%�I���v��X��
Y䅠|c/����� A��UzRIlkC��ؕ�5�_>'�7�I&c��:k��̀��s�dk��)��hrB��wVgBy�ϑo�ݠy���xe�!0.��K��_~� q���x����ɘ���a:i�}�Ѥ�#�YЫ>Kc��}s�ˋ��1#I�M��H��ހ���Duh��LLIV�Υy���{���(�-"=l5��U,��Uv� u��9�>ڶ P�;yM��D8�8u)�䱹_k�>L�M�k[����p�U��l4�s���=@%�����}��-�}UE�!�,5h�Y�z����)ܱ���C8���I�mrE��B��KP���`}��=��,psSN���劏)p|��i����4ꃫ�V\G�88]�^n�[�{��G
<�x+v�x����W��8[Jy�;h�� m�ŷQ[�U�kg���4�f�W}l3�K9���j�Y��ˢF?���V�A��~P�C�݇�X�i����IB�_[o?R���n�5MB37}����zcmQi�Q�%���wZɣq�'�����	z�P�,��}y68j�z�aR��"V���I���j}po�>�Q��Z���{`|S�B�������
��F�B�|c��nE ����cԪM����'�����LsO3�s5�(3{���	o�D�'�B5��=?1��X���T��-h��僇����\��!�AJ�,_ ��FK��.������Y�zݴ�����9u� ��~u^��-
n<��}%�>����u� ]�n�Έ2��(��]�p5f�]\��Ѥ���I3�ѿ$>�{Vy]��)��x�̮-�����
mŔm#����Y�"��2>2���g��╍�j���t�vJ1|i�@�P��]��6��O�2���4�m>�ʂȀ��=w�N�ǅo�rCs��)x4���M{�?�=���CU��\<�rd�-�=	qٱ��7��f����0'r��@�N�N]�t�Ƚ��,�6�����<��4#W��ى��5Л2�O�E�𮣫��%��������s"3
�6��6��Ib�����^ �q
W�+؆���&�MKU��v��(
�:Jլʒ����?w�}�FQW��Vf}l��ԿC�u�T\{��5��Eb�Ȁ��f+}�s�l!ݜ7=���8�4\4�ե|v��������b��8C~�娌��$�߈�w�>+B� �
-kreޣ�Ѭ�Ɨ�p���tg��r���f.&jf����C�9�*�d���W�D��#���Hg"�A�H�tZ�>�Ma#Xd2��o~�K�nWKϏx�*&>�,n�mG��f�����tg�����,��b���h�ɠ{�MZ�w9�ӹ8���u���3h�����eid��������_IZ��	�s��!k���sJ��IҎ�6tD-��E������s�W��ZcO�'y�qF��~ûl�@��.��3�#�@	������1c�uP�ϱ�����9��O��f�>�G�	"6����w6꼶�l�HQ��� �4y�_�����m1�K�i9�l�k��	Y� ��>GƏ^G��)A!_��˲�<��!ӓ�R/��F�\pjTdؿ�0[�P� 3 *��ߗ�`�n�$�gU� �ｪ���Ll��&�8��2 �]�zɽ)���.�p��V�ݑ�� !�}K���"�o_/�ͤ�Z� ��:�$�3����z@�����r6m��ʢ�����f����B������6�����'�j�2��?l!�+��o/������J������V�;�L�Uw]}G�S�'��q��u��^��w��j��||H�*� y+�;�V�B�P3 �.��{6JQD�OD���;E�<��a��H�*q�l�h�����%eM�s c�~�:�}�~r���%��b4b�\\S��M�3�k@�o�h��q��y�m��_��W|y�g^'k��I��pIG�L�#G�� ~A������z��O�( �zʑ^o�Ꚓ�\��b��t[ �d]I�V��?����ݗ��u��O6M���5 ��ibݨ��j?ha��ޅ����2�hyP�A;5�q ^����N*���Fc)�,��ޭ�Y��T���M��9 �T9v2��"gG��������8�ծx�*v,*�/j�c�|Pep�U�����6�,Xg�Ew�C�r��t�O���b�Ĺe�u��l� �j��si���g����u�}w��d�5b��
Z��8|��ڽ�ڦ¶������v7�-���1���'5��Jsm6�`Szw.�5 �u��r�?�Y��-pJ�k�HLv�s@�ŕw9!E��9O0tN�����o!���{��6߷N�쏅~��i��b
��NK`�k�9�,����V&_J�"C	�֬�t�Vg��d��@WE�O��>b��E��&�����.K:��&�Fu���( p��Hoa����&�P�W��FU������k_�|1�!���Ϳj�ʼ���ÔO:�CO�YU��0��0P�j8 �|6n�=���">I@�/+D�_	3�2��Y!$�����3���u��2#ڏ"��-cq�YȆCF��:�f���;&�y%_�W4���&������ş��^vC��F;)8	G�+�d�Ja^M����`4^��#J���Z��я<�(ìn�H� �{�ep�$P�D�ʲ������N���ܵ��ܙ�g��2jL���Y�
����o��;��ާ`AQ{l�'�,	R0�P�D^-���Ɇ�^�%P�"�l�����ڦͿ$�x�M�'�X�wi��D�4��.�Ď8 �)�	��kc�����T+��2�ۨ��Ə$w���5Xww]�����d1C�"L�J|�f*qw�*�1��zZY���O����J�i�PщԻ"_#�Z�I�S��n˽�Q���`�Rc*�2��)�}�2CA��W�Q��a��w
5����77tRM�j��'��S���B_4J���%Q9��2�[�@��B��a �*rQ��5./)���F��0�?�(�}*�L�Y��\6��.P.��,��z�C��(�B tY�Ex���w h�j�VFO>(�#EӜ>W�a������� 3�S�:w2E�{��Vg�[�Ƿ���9уz^�pOx�ݵ&��4|,k�hշ7�_ǜ(�T�%{R����X'#Z�R9�b.7�L����+��64�7QA�'��IG�!ip}0=��u�*z*^5D �8��&E\)�u�Q9|�<�ĕ8Y�(�Y.�Rձ��|&����~�� ���(s�(ei ��Ԕ_G�,�{N1͡Ӂd�aݼ��>�X��u�Ւ�A�ZN��� �죥A gjd�'�)�����蝗��Ǭ��a�f��$X���;Lǵ�/m�b��t"��q�{�
�d�^���s�=��`��k���Ӯ��^w ����N;�������/DX��z�c�����P�0iz�����Sl�8E^��!�|+��Bn��"@we��<�l�0$�������2W�5"��p���������ś�ƃ=�����x��/'Yx�`wǚ!�t�}vg�j�7�����e�d��)�`��S��XmP��z?�bVԙ����(P��7ԍ8����ܫ1�S�%0÷�K]�K3x5����=�˚L�;a���Qclug#d/#�O�p7�,�@�����8�<$Y���\9)A��(���q�����鏄'@��u�` ����8~q
��O ��Iy�ewV�����h��킲�'	�e�)�՛�.dI�Ҙ�v8Ó]2��!�8a&��?~s;��pJ�-5�Â�&gRW�¸��k�v	�+",�1Qz�ׇ<���U�X[�I}�K��T�5^E�e��ԹÅ�y����DA�!�>
��~a�lW�h5���?���)�$C�Nȏ���6V%�D�B�{���VC#/{b#�>���V',��v-����[��X��9n���Je?��B�7q@�aM.��Ŝ�
z�ذ2��zz��"[�;%�Ղ;��zCz�˺>���r��%i�=�&��8�ڪ�Q�ˑ/�.;��&��0���燐_Q ��j��9�C���жU�,�=���"��:��p�Y�tg���"�*��L�[��w�6���R�c�D)�l� �"�S���>�ҩ������VDD������ǥ��f;�$��Ie��"�䢟"+�yr?y���y)aF]=0��B.c '��ϫ�-#�j�$2d
��ZM�F�q�|ϸ�����Rũ6��H˯;��}"^ٔ�v�N��fݹ"�y��쁳�U*��{	�+X���>͊� �3�_a_�����y��:b�oy�WVv�_� h\�@���0�&��F�~�E����T��6�(0vKb��̋|"�����8t`�r�h��fFbC��Չ(�Rj�y�^�����1��
�24ڛ��ؙB4������2�ĺ�nu�~�B�=Y���!sΑ�!��b`'L�c؂2�����2�R�4�κ�#�S����@g]�D]��3�@ֳ�%C�j��!��sTq��]J�k8n�[4,�ɸ��K�<�e �7�O�OJ]Q��O��AG�m�Pʝ}�x��u������>�A���ݽ���d~��)e�#�z��}��d|��JH�Z�6P��Zg��̶~#{vłƁK�po���J��P�` �u��9���z�#��4��� �K���K�� j���U�p���B$|�����%�����h�ͳ�R^�����](����?���i���R�<G֥�M��<z���j�ߑ��p�ݚ��Tٷ��b��~~��'�|��м"a}�{��WE��x�����9<d�o��)���r" ���W�X�w�Mx$��C�e�Q_��0�`�i�nº*-s��)X�*u�]f_�Ow+4XӞE!��9p�`E����=�ɛ�#��u0},3a4B��N4��v|3F�X�3��������}���K\��Pkl���X�RW� �k��b �r;������p�1X�B�m
y����/��i8C��c�^8�*ľ�Ԕ ���Gr�m��.�w��I�ܬ��s|��=�h����QH/l�UCM������_�c��w$�+>H�=��n�poj5Gv�Aє��sR�
0D�c��3��=�SN�B��Rv�q*�ju��)�݉��7j���g%4PFZd<1�������}2��s3$� Mp�ݟ\�����枪��C��aۯ/+�kL�5dt��u�&[\���cb��� jV�S�x�PX[y5V�/�%2J0�^4����Ɋ���V�{}r�ϩ�(J�)���qm�����j?))5������92%I\~Lřc���љ�o���RK@.���&<����?����K=Z�F���ut۩P�����b_r�q/�E��7`ch��
^ʚu����Y�,D\��܆��	�ȯ�俯k_2��ߞ����v9�y��js��nuF� �$%O�$��0��ﺖ�� �ҽY
mc��;^�~d��	�A3��6�:����@mn��듼u�� ^6���fb�ԗO}��1�Nu���ڣ��e@���.'�또����ݞ�f���[3��vB��'�����0��Gi*n��2���
��q�J�pS�8&�����	�]��_'���b��z�b���[�'49U`�L�؁lQן#�v��}��>��9s�;Y1"�ڏ�lO��#s8�ت��"�����0�W�b~ϔ��E ,�[������U��(>�*�,��h�)�jx	0����'����5U��hg��#�(�'9�w�gq�'X�^z��2��l5Q�ާ�5���h44�F�yV0�۱�9R�)Q��T��l�B"���?�)�˙;�KVÈRC���X��'מ���T�FN�-W��K��r�T�*���58�k��mmM��[1i0C+3�)1�h%P._7���d�AT�a�K��˨����P�)t����d$�茯x�Ù1���F�A�B�h*�[!�& v�N�.����� ;�!�d���2����?�V��9nYh��4�Q���1e��v/ nrW1b'��Dp�I���G��t-BL3e2	#�*�����H.CO�`�X�W!8:�����\�jlx��(��xh�X.�<h�)����?�cW��� H�o��:�π������)$v�k�.^NDZS�x5I�>y��KM�����7�����<�{z����Ŭi�(Z�EG���1�AH%*��]�NB&�|�q�4j�~��W���#�'pT�w_�^|*r}��?Y�'d� jQ5�@��ޏ�֌���//g���\L[���Ġ��D|���\�\4'j �i����E��ztN?ԓ��u�j��x�G�ȧ&d�c�|Y��Ce1K�~�V����U�R�)��+e����������>�ĖhX���ʏ�x���{A_婰��xucƻ�)�D@b�����(vGfߤ��~~�ӈrw3`/�X����F8DZO�)�5x�6yIs���-��/'�5��8�<'x.�)�ۄ=�UG0���[�	?��i���~�<�� � <��nc�kdk���v�slѠb��Tɘ]���S�>�q�9���a�W�	�s�&1�1��C�� T��7u?@�_�B��&�̬l�T���-���ez**��o 'm1���-s�+8��M�u1!��	nKm�b�[pט�
K���f��{��&��w���4:��5#�M�FH��r9V��Θί����f
6�ᡧ[��C$�U��U��J�?�����>S7V�(k=���Z�Ps"�}g�Є�m;��S�R��	���l�M嘤H\�=�t.T��FmЭpG�պÔC��I�: ��ޗG,/X�ƕ@,�9�n�^���]���=�AcQr��b_
$�킶}mLe��+7�ܰ!���v���7�K��r�w��xj�
m!:�N�i���|�Xݣ��;� ,
���\7w��-a�\[��d!$����cI<�J}��P����w�D5�;>�N�"W��^��F�p=<�Ǒ!*�b�k��������R�p���Ԥ�����|����B�ܧ�dng���\���-���r�~1f@���y0�D�LF���gC<����{�%f�j��^��-/��;�ʐ'�s�ȗ��J�lH�!�K
�����D�o�G�ٜ�{��{B�IM�|����V�)\�3��ub�b����|�^��d��Ԟ��5j�B���ՁH�>��R��Ck�{�h���2?5��m`���x���G�/Ӈ�S���Ut}��2���Wp��h������������ws6n'����g	$���\|����%�ƛ�O���Hw@�ϐ��w���%6�',�D}Go&	�t�	��J����#47H�ʌ�r4���`��tWL�,�����D�8���3n?BO<���	{H�4�e�rGG Ya��?�gqS���@�sW��ł%��O�%AEY+��~;���ń�T�!;�������I�A�x�κ)����+N|���!���^�ql�>*��i z�eqB�|�:m��zh�;׍P�͸O' �V�K���h&)n���mF$���Qs>�p����m���mgm�cYz�~��4�_������d�6if����x�"Eb�&M���N����NC����$�ŉ�e/�|��CH��6C�K�wc��d���ԏɀ��@��h�݄#B�ŧPjk<^z��g�C��>#@��{�Y:ļ/��(2��R[ }^.XJ0��'
ؿ��1o@/���	:���
�^�EQ~_�:U�m�����ݳEDd�d��XЋ6���m
j�e^�鞬���%<Y����Z�R�+C̭_ƽ�|02c)������gH�Y��m�bO�p��(x�:4�A�0Ɉ�h�Qr�n�C�ѻ�OPn��LHV�� �{�6�M�(=7�S�T��-�R~�+�ي��?�+��<Lëގ@C��{-5�����O$plEpG/є�#��&��1�o�[di�e�(�اv��S
��K�p�A	���ʃ���;�?���/�H�'�$������{��S�1�hh�a���bOa�i�	�7���#}�4=�������}V�~�J��g���S���.P������'m$;+LZH�ڢg��\�k��R$��H�T%���y�W� � �Q+���"�F]�K<�&n��9���gr��2<�u{�y�)�)^ ���d���-J�Fz��f��z�s�i���T��mH�~%ʡ��D�����7����!V�vC�� ��f�mNF�4�e~�\��@�^7�ͭ� M�A�G�k8�UHNP!ٷ���-8+��o�{�k��'$�j����,K"��ϥ{v��u�]t#.�&���tt~B.�s3ю�	�
�Ki��4�Gy���>�����N������ ho�C�i�=|d6���U':e��r팢4��T�ě�.��x�Sh`���msJꝿT���F�YtDk��t��R��Ux�����P��V���S�;�SsF<b���Í˂a��H�j�	:s�4����L����@Y?�a��k�n�	�G0z��OP��{"��KQ�UUv��c5��YD=f�� ��Qb<�W�1�7*�]x"�y��κP <����Ȝ�oP�>и<�xJ[��t��5�Om�r��P��RF��5�ߩw/�j׼�A�#>�;�K����U�TJ%Jxg��~�ol�����3|�}?>{��P^�R��V'�����e_(�����}	�"���LF&�r�-�o��j9g�������c>�ŰK�I�u���'9������J���b�՛Ҥ|/^���t7hE$=\2V��SꐸQ��6��	A��y kL	2} q����D��[���S��n)�n)J����I��UUn� 2�N����mlM�7�ܐX%ŕI���H��^����������	s�u�oWF�ZUp�������~����d�B߾煬h�S��a
�O����髆;�S�������0���{D#����њp!H�f��\�H=NC�<�Ͷ� 4܋Nw�q�#��l���y��7�3�44q�f�����4T��~) ���F?�#�K*����jn�<�\��٣��� ��G��^�G�9��;y��6E�&9\��*�(�=b��{���?Q9`g� Upv��*<`)v\$��Y�����.��62��-
�? }2_f�u�����0�#oJ�ZYfX�����|Sy�M)���)�g����	�����9� ݜ�-~�ʳ]�'�����@�U4�J���T���7V�wmuv�0Ns�§t�rBqӲH�Q۫,l��^D��H>C�r�a-Р�/!�������j#�0�W�kUrqd���׶~�����z��CK*��g�Ub��[~���q��f��eFb�
�Ry3�#��2�4���^EKh�V6r(Gć+�h߫F�w��.��/�O�o�^,~�C�B�?h���[��UR�V*�8���l��-��ʻ�yZ�-�?Yw�?yx�}܁b�xPRw�vT����8X"���)F�bo����.ʩ��n��d�(�Κ�S%���ٍ��)#?{a�o<q;vZmg�i-�ѳ։��j� p����/|b�uL}���aX����d�}�D�������x;:��j_�Q�O�����5 ɣ��s�Q��W����4�cr�5��>��<a�9��t�c��x�e�Q'��&)(ۅ�mr��;�������k��1	|����r��c�H���^�����vZ��2�������V ��a}8+�}�(Xq\�62PR�6p�\"�� ��`����i��>7J�
~5e�	P�!\�ө��{�\�����g 4
�{�=/N���y�'�j���p��˽�?&o�5-_m�V��V�����5!$U�)5�kR����X��k��C�A�7�x��N/�'�����i��i��(����A]��ҎH~��&�{�;�>Ob$&�{�O(SŒ�h
�0'g�b_�� �����4�^���H������
H�D�#�2E��
E<�vR�\39.ﭛ��=�*������K�J+���M!��,�IhPN&F5ϋ�bC��L��˭�-YϬH� �m��6�W֓~T��ׄ*�()�D�Zh��s�;���F��q���*�W�m�S&�İ=OK�&�
=�� �t�0A��"��������0y�^�`b��x��^lP�(ɫ�	��$V�׬�B$ɞ�ؔDߩMF`3NN�F�ZyT�� ]�y�K�M<�[єT���~��J���pHW,⍡o��� �Wq���	KJ^.�F�HЩȪ��Y����d�ۥݹ��E�*!�;#<�}��A��r��>4-'��\\,�\Y�u�źJ���7�_䮩��a�y��H-��HH�TS~Oz�g��E�8"j7T�
:��,��*^)Zw���3?��4�J�7��q�:o7�����Fڅ��3����+rޗ���[k�\�e�;j�S��&h�Gu𑺈B��i�ْs�(��O�N�aF�ˁvC�D'pL��I��grW��z��	PԂ����C�4�0����~�j��	'R��r�Q/��݉�evB��0����}�Dӯ�����t͂�g��w�]���<��6���0��>.�Bx֭a�Th�	��XIi�1 u��٪0����El�u��k�u��?�]�*H U��Թ������sH���M(�3:ٙJ�8aX����I�[zgq�K�i�J���OD�g�����K���HW����=��	76p��e�xjk���L�G�Q���"_������E�����p��B�A����y�t.�W5�8�6�l��è�Fr*Ls�+~���(,���lj�3�^i�_.�4`iV����W�e�����}9�z=�(��l����x��y,a~�{���˶��3r� �2�����J|6��,a`����:HS��ǭ|��E�<��B�f�**��z]%��s�k�gA��p�RVM���1�d|1�:5?�Z�C�ӌ������c&f�m�L�O�/LE�y�\,|%3Uw�U�_��t�g�Ե�g�]��R]�g?�t�4C
�8�U�~�2T�33:u�/u^p�4 H9�l��M6;~g����x�ză{W�I�.)͒u��8�~��7�?�>1~%����R�"�K���4�m��-�ϡ��bN�������������@*~�t��'�'������x���v�����;{x��.U�~<Z[�ee����W�̝=�L��H~R<�oL������P�d�A�D�#�3
C0���5r�u�J6�M��X �ni��	���_����ƽ8�[���=G[m���?�P0�g@�&Lf�G4�3)���8>�/��G
~�&�]X�]���;���2:��K� R[� y�OW�m#4����@@[H�?�>\���,WOc�>�%�6[Y�g�k\|C��v�3��S� ��9��d��?u��ҔAJ�YY�M��},��KE�UIP��Ew���N�=`���s�ȴɅ;c�{kݳ�}X�5E�NUv�-4��{Z�̆����g.☿�5t�mn&�x�!�E~�\G�m��@ ��ȷ��Ôפ�{r���T|���ؽ^㙐���=C�;h�6�H���~�W^K."��D/07f
�3н��d�iR�GV-2p!�,��8������"���{���X���1�xvR��*)���5*����pss�H �-�_�|�F�\�똀�j
c� ���� :}����}�0�;��a��e��p3I�-2�.��D���c`�(�3�MmDg9��R��~Z
�fN2��8�����k.ma�hF=3b�c}m¡%/�Q}�����q!ř�ɯ�{�!*�ڧg��')4�{��gUS�BbJ�d��L7�H�������C/ʯ�܎�}�e��G�����
8���prB��Y5 �Dc"��}���s�]�P��Ȑ��\�k��(�I���m�Uh�!�f��M-�GbJw�̤��(J�ߘՉ��ʿ�or�ġ_}�}L��|���q������,���C�y	A许'��d�Hw��>�S�dq���<�VՁ0�&�H��ÂN4/t�wS�.n������k�}�xw��{jC�l	5�w塞�0�ý�d6�T�s�I��X}{�˂k�¦�c�cA�')�ZP��u���2�%=�� �h�1x�'gޜ�(D	o�q-I'�W�-=0J],����A��Z�}%$��m��f����[��%��h�M��F@G�CŻ���5J��꧳NhU�7S��4�s�g2u/c�&F�^���6S����:�!~V� �;��r J��Ux�Dwc��E�T|	����#�3@�<�*�k�$��Q
�����@)���!��J��˴h�=%x��MC��0ǭ�8�G�	VqhP9Ɔ��;�3�W��#��5������`���4z�	�����̹��ߍP��Y2��� V }�<E��K_�� G��k"�Mlq�-�{L^Ւ�->@ޏs8�FW�;7�	�C�y�"��RM�>q���b׆�����rPj�<��h&ar?�zDU"[�#�t<��h�UUVV��^��6�n_��,f�,ۤ?)w<��������BQuz/[KѢ�|�K�Y+
���S���T�iW�2���� ��dik�;�{�����0��V�j�$3�)fN�XW�3�p�	�	q	 ��A�J|~
�6c�»�H�$��dz��/�75����E�t�Yq�Q(�s@�c]��.mӴ�5�d?W HA5�&�W��Gn�m��%P ���M�(�:����Z*��1&�6�P��-�6��*})�� u,��H,�����N"Q����Kɞ�Z@7@��ϗ���:R/�T��J�ڸ�X�����\b�vWF�O���k�����|i9��J'����r4���R�,&��&�Np<���Է��P�@^�Rȑ�@�ufh�)��T��]Sp�p��(��$���w�M�R�L6*Q����kHo ���Ua��J^�*�-
J~�]�3ǉ�&c��y�C1L����ږԭ$��)�8�@��;y�H��Wly����*k{�U�x�F��J@P���w�[��3"+�k��1s��6��듹ū�O��_hx�E��P�����������v��J,�@�5�9��a� �tp�@�b�u-��Xт%�ǔ�g/"��dE�X��\V!-��ܶ����EymTN����ړ�`�.�X��8`�����>�-� Dyg���֤���OS%ݿU��!O���𴙧s�H�^�rg��� /���o.����5���g%�Oj�J��6��$����Ux�dO�.J9)�A��$<�V$�eP�$�#�=�Mˊ�c���Bu��U&�~^F���ȏ}�\�Yn�l�P�{��
T�"M5������y�~������d�}�	'AR��mX�*�2ކ�I�1�[O�-g4�
|�2�z�846�5���L
/S���V��On��K�?q߭�EQ�q��n<k�Dw'�N������djr�!�q�{e�F5?��+~/�ـ�>������U��T�� �['{�z�z���Q��em�e�4o�)H&5�J���%�$���&V�5�[��"-ݧcw����$�A�-�_�[+N�r��8�_�������;@e��C�نh���o�$��ٻW�-��-�(W��4X�UXQhI�nn�3"�.��uMև� �B'��K^�Y:���-��X��� �hEpml}p�:������VSP*ѻ�}�:۲���*�~�}�gH@���/�i�=��c�g�;3��*YD�ՉZ��I��؁���TP�L�pQ���R�'*O�U{�C��]+��PF��M��P���R��5������E�G�gvhZ�U����s"�Y�<��Z����ژ��X��ߕd��m�N ��x�y�����#�����['M��B01\ޟO��Iɦ�j����sj6-�^������5D���͓����_�B+c3��=W�|C�Y��(�Qc�l����f���\W�����d&�^S���Im��6>���\�1i�ѧ��:J%�^"�4�B8�!C@kۢ|,�P���w�:s������^5���*�|�1`���Pl62���G����W�(v=��O���W�tJ��Q��[�TC��u>A���`��ڋ�z�LA�7��(�Dw���N��F+���bo4q�s)%u���t�����~�J�E
�������R���<������0[�/%h��u�/₁�'�Ċ��<���ݤ��D�����%B�l}�e��х~�t^����qo&~��"K����E`cU`�)�'�u�[��C���>�6G-^j,B�h9�iC��Ӳ��9߄>�M��l�V
����j������1=���`"|�r{R�5y��w8�H`'�����[���ݙ/1a�3#�ʳC��~���"�ݿ�-S��=���b2�U>r#>R����l�#5
����N�;��z�R�_-9f$�m��L���/o�"|p�`��2qk��l$Y4�j����.C?���9�������������oө]1�@k�>7gs����U�k���tچHh���	u�>��Ax��w`�Q[t��U��,_��?��ʟN���8�SK������H����7(��?>�$@�����޽�<>>�X����AY1WQ�s:
nc8۔��D�c$e�l+�|�2�C�ڨ_^�$Hpƺ���'�l�Uh|��&�@����&�R����?=������A�OD�k�������4�K�Քe�l����5����1b?a��L~ZY!,��������J��<� ���V�g�f~6�{��������
��_U�§+`�9�\6�p���b ��t
� l��L��G�����	��@�ka`_��ec�Ո��9�$�Q8���$3���ޠ�לۍ�����Eȡ�7U���}���;j�� �3#��0��2����ű��y� t |�|.��]��%�>`�N���a���5���=�	5�'H�� ��R8ęPWQ8rk�_WCH��R�2���^�5�b��j�j ����#��k�5�gN�"c3}2+TcT�ȵLU9bx�y(_��TK�!���	q��|������I�XJ0�<�f?ט�g��B3o��g�k��ȩ��d��}=5�6���綏�S���F�`Y�?g��Fb�`
�.X��2�8Iс�Y����+\zl�Y�~n@�o�$dV�<f�B��%О^T��a[��-e��A#����MW�_8��O���{���'�N��ew���?~_��=�m��]gO=ު�3���QED$^�݈UH�1���#�_�=�d�ĝ�![N�,s�����ݣ%�*�<rv���̶�t��TX�s~�`ڍK'�;�9��Yg���4�mQ���C�&!UGt��z�~I�E���DLMFvR-za�ME�(r����c�_ 5�h�D��4[1�0�Ҽ?9{.y�S��)�th�/R.���=$^�9�M�����F��WS��R�ل��Y\�6߽K�l�ixcU�O�϶�W��Tr���!��>�0͒������2p�b��'=���}y��l���5W���+d!p̈��R���JY�{^����"����Z�6|���Q�or�T�o;�r��(�(9v[j�`���1>Np��-���$�ێ�s����,���g_k$���&����k�.�Y��.�r��O�6B���q��:<��=�.��s���t���m��@��K�.{��1+HO�1�nH�=�0I� �Ҏ�C���,�V��6�u�� ��S ���o�ު��7
_��J��^��/������̵�~��7�h�YbM���ԥ]d(��9eh�x~��e�yr��g;5�G���ok&^P ��`�#m2��J�U*�D�c��[T���@w�eeu�3�
}:�r��,�lo�2���U��]:�	�V�;C�	僱y��m�Ѹ8�_��L�M��<V�Y���p9�EZ�%`��%���b{f�.9���D��@r]�m R9���SQ��G��y�X��^�-���nW=U/�������]LL徔̻v�`ؐ�N�s�-e�t�6(�	:��S3�5/��s�կ���66��o+E,�uS � g��H0���NB+ŗ�q�2�#ۍ9��3&��Y�*N�ZM!C��)��ى��-pL���b�)@{�7�"B�,ṓ�3�_?V�ȧ/5b�����b��f+�9ӓ��{�xϜ��wbKZqΘ��� 	�hM�o���޵���TU	j�:Ѝ!����+IM&6+z��T������a2H �]J`�]�+H+21����b-ImJ7��POf�p��{���Ϳ--�^.[Y3M���R���mT;Ye�o�i��S&"����Ab���TsQ��Y�]��9>����9��+���~ �H���J�Չ�b�c�փ����!LV��WՅ���hRj����-�O#�d�wmo��}v�
�YgH�R���(�F��xmE���V1E+���*Z���W���S����n*evWA��]�I���I�{�U���q([{b��m�'������>`ɉ��%sZ
�|:��B�ez7u{���\�P�gNm!�ԃ�������G�Ѵ�qӀ���ri�kx���\�@�d˺�ƪsg��
���]5�C���� ��\�ά�\���P:�3��T(?��5 �Z�Y��8�OG`��Fa�ra9re�킺*���̾�����{�F�*�Ȍ�j��Ox��M��{b��>d�Pxkz��+���$�ȓ	"JS��i3��~���g-��N�6�f�i)�^�%Y>q´%bw��t��
����ķ��S�p��:(
�M�*���$0�Gп�Z�Z5n~����}���cP�j�Y�������@����4�
���S�J$g]F\��뺄{��M�G	@��=6@���۪ .-�<�؀���� 8ޫ�3Kφ3��ӗ�l�IƑs��Oʆ�n����y����'(�B���%��j��v����#ĭ�G���+��wז��ry�63/b˩�R
���K�nV��F�Sn��O%{Z�x%c��r���!����_�)b7 0����avs��������4y�K�+8L[��������ZϐȐ�9x�~T�KV�k�{�+��_&�cQ�uP����U��0�J����Mq��n�	�x]����*�^t�Me�����|tN��&��,`|6�sNTwh��|��N�}�,�?����{�KY�ey2���Ì��R��9����'W��MKRZ�������~�Ѭ�������Z���gwf��R���F��מ���s��)�^.��%���'��W��|P��q@�8���f�jA��zvs�FQ[T��--Hut�\��4��N`�SaP�~��@�E�v�B�:���	n�b�l/q���2a.P}�� (�I8�7!�H��i+���ԉ���Q�z��O��t0%%�]���^��kVQ��G4�*�5��a��䱻DS��J�u��e��R�(YM"�ױH���
��<���N����.�?�4z���@	��h�¢��bҤ��mgU� ��ｽPB��ȴڟ�p�QZo�	*`��u�?�_�s��Yrt�I�ikY˃kzW��C�MI���E�N�4���:�����CV�1�K�/yN���'Q���$�0�"���b�jz� �:���x�3�[�6���M�K`�%����&��kX}P#8�R+�/�e͘#1ڰ������b6C,G��f�=�9�G t���t��N�����/G{I^���u��s�2��w�W�����>� O �H����l�.u���>;��`�T+4��g�����0�\�g��ӽyаA����;�"��n���U��v4�D�OO _����<yT�`ը|P�w\
���b��a<ڤl����@�y��JQn5a�bx�Y2䶑:Ӳr�����D8����jK�����8x�^�=�ͥ�WŲ��a�����?�W��3��������k�=�Pe^zQ�ϧ;�������ڇ��[�m�ɰN5����Y8LT������~{���h�qd�ì$�mj�P!��]��1R�")0�ٳ�滒J/|�����TT@��i�,r��*LN]�h��e���=|z�r�������7����	%9�酏�O�Ur��+��,𤿮l��;/*���!�8E��S�~�1��n�|W��%(��'�ܣb�-�=!3�m� ���t>�͏bWXQ��Tu�p�ӎ]�ˢQt��E��Dl�2��'������~�x�'S��ݰZ�r�ͻ�]i嬝h�!�����=�A�O���,��Gbj�-�#�SF���S��9���Վeb~u/oM5;�v���_�K��S��Q,����"�E�S�5����4^�oH����
�wX�*�=�1���S!bj�W�h�K��z�=�g�C!�9�	x�Uԏ�࿚�t%qC�me[j�K����*���?���]����,�JA�]6��e��U��fq����E�*j�vm�B�B��(j�����b�ؓZz�V&{�9M�tF�&K^t���D��W��SL`�/�A�lW��X�	+{$�g�ò�ٷp�*�._�ɉ%�Α��������������w�[�8aڅ �����4<ZF�J�!��x}l�r�y��A��4�����&�rl��1�9���nFEÎ�1��3)S�Lg��O�������BR�,R_�ˋ�^����Co���X� HX���,�&���k�~N���V9��8���r[o��v�m5��P"�۳h`���oLE�L���D�>ojF�Ml�a���qx���.�,4K�O��s�u��^�MN�g�A0O^�:�7=%R�L�-��B�"���?�;;β��s~�78O�:1/� ��������(�x������'u%��]_T�RW���yk0Ɣ�����@���_｣��%�6$<�-��/���b��Ȱ�����xX����K^	)�聚�4?K壚Q�O�+ez)3�ѳ y����e�v�wњ:����h4������*;{���,s����ϮEL�yXC�w_Hj���a��:�Ϭ�&Z�P��ͦ�2�}Zm�&8V�� �ly�\��E��nm��U^�D��ai���q��,�i�Y!����
�w�h7�a�d7u+ �C�T�VP+D�L���bmDΗ"�nr���SXU���X��v��W.L��Yy�5.�<�L�x��nx�;�c�I#��*������\�+^������v��r��(����
�M��'{U��u:��:>�?zO���2\�|IQ�BE�]#kf�u���a~����y'�49��-��#(� d����������E�K��A�����䦊���[��Y2�Y�#(���U�W��}�v��8�o^1�e���-wq�[ � =�*�@�U�f��c�}A��ɏ��Ѓ�7a�-%v ����@Q��<~�����%��${Ur�O��(<:ޝ���	�\X8ߍv��]$���H#�Q�+�N&o�뾁N���.��y1s(����6$شD�#p�.}	VП	x�#ǹL�l��#��*"M���i��=��ҫ�`b�*��8�wEP�,B6)��R�w�l�|$j ڦ�㭔�#�E:hED+�/���̯� �am/BO7�J�nE�`y�3��F��?���W��0q�'��O�������v��դe��[������^"O
��z��1�ok ���$Ul�*0��I�F:f`�tW�+���֡�Ң�6����5W�J���y�P���a��Oh�k�Ь�q���"7y�؎i#*��4ؾi�쥏�fջ�er���36�'�hr���_�1��b�4� ����_�a�����pg��PЧv�\�е��S��=��*�ׄ�s��� G+E��f��!We���Wj���%O�}����8��DН��~2�jp�X0w�V�����<��AF�0��/��� t�] ��r��P4Y�I�f=�ΐH��sο،J�����0�]�&�ш�]�ϰ�
��020�.����
+�4���A�<*bh$x\�7zS9�,�i�SƇ��n7LU�ߺ��NE�'��Vl�VD�����;�!h�c5 /N�8Bl|pQHp�˸s���Q����x��ݧ@�} ��1�5}E�+),k��2���4¸v����	ݠ�'~�Z!���ag#��8�T�݅I����C4�XN�i&���:�{bf����<%wK�T5m���Ç�[U��0,s6]��N/������r�zTHP�[R��}j/�q��������4�?���g�b52�T4F�.��؛g�=�]/a����ؿ�8�L�6w���nDAI���3��� "�|n5�{F��X�e6�E�'����X�c@�� T�?ښ ��A��y�W^�'����B�"*lN^nh~}���y8�]��>]��g�<6Ad2%h�?Q?	̷��b]���8?C'k<�#�!!D ������hj�;�����,G���u�{$\�<qZ'��&ND�p�=0��y>"%ޙ/)�����w���b�������Q������eWT2���?m� |~�E��;*�ŇvK{|7[E$q�9�|!	A�KX����]���"nD��ܴ7�L�ef�������{�CH,
�����1\�7����3�d�)���\C>&d�FTb��j^������k$�j�vg�u&Ri�Cbh$�T��,�Q$�9�����hL��񁽐>+�.,����4���jB���m��_W��Z��5bw� ^�`�Ճ����;a��rM�TdS~t�·�wG�QuN�E9��8�%�Փ��n��I�rx��s��'����	>,k�0�w��MHtV��F\��T�b۽�$Q��W~7㻱��u_�Dr����"�J(��g����� ����a�g�g�fx2j��^���GJa��T�T��A?�Gb]�����W�X_=bSȍkB���&E��E[�$��j�ѹB��ʣ�� :#����.�Y�|*Ye|}���J����aZ�ֹ��I�%/p�uR�k1�4��8��쳙���.�<��}�ˮW�K���5��d.�9���Ǹ6���J�)b6���.�Y��f�;G�u�Ҏ0����6��ԇ�������^�+µ@�]6�*�4R�p�"���i������o'� 0��x�- Խ��Tjx��"rx�;��8 �:&�����JZ-�rZ���*��8~�6?�S�3Rƣ�[z#x�m�n��h��1Y@�J`|�qI�OO�xd��wV
Y���1]N����Bp���r?赩e��a���IO������˖Q�B��W�;�UQsv9��zF������E�R��]�F�x���~,^��X�§���	���^��ݷ��XQ�$8�$䥒h5�C�]���y=�Z�i"����L]�\Ycة=��Շ4�)̉#�3uf����lU�f,�&��W̆�9Px�ܨ��hؙ��`P�a}�@��A��������|t�)�Y�}l�c�D|h��)���a��\#�b0b0p\ȽpnO���������L�M�O�#��ۯ��*]
��[����h�<��v \�j~o�vy3�\��	����C��v��N�UCҗ]��=��xKR�;}���<������4�V5Y�-��O�z���*���3{Jp�ޙ���b��Y*1e��g�E�)���[���0J�.���O0Ǆd��)�q_�$�[����D@��3Ū�/�PY�ï<W��U��Ш�><bY���6������d��P������OW���ٟ��^�b�X���<,R�7?T�W���e$W�0�~��SN�co(�p�wXp��J��5��g1=}�H��9\/'Mݒ��:��J���l��(���(�m�/� {���=�H�^!U�XLhvŕcD���`dS����R!�~��ȧ�%E��Ͻ#��v��8�E�Y%�mP�8왙����m	�ra���-g������x��Y![�!�f�������ٖ�A�mz�[H� �k��D�5k�m�����^N��+2�Pn�K4�1tt �f'��q�r'�j[�+������b����4p�ӱ��åk�� z�W�%��D9a&?�}��*�bD&���OC�Y��C}�p;���w��_�۸�����j6o^jc�Z�
��d���A�6���`տw�1Vl�4`K����L��o5�},�j�]�T$:�C&�~�G�b6CKf�N�_�}�;VǱ��Dw��f��E���@�^����g�}aF�i�p�4۪�՘�"�mOL
�_�:��9 �{���3�F�c�HgJ�TS��5�EPC6�nt�WZo��ʋ=cZFp���(t�fu�%�<���q���e�Qeص�1T�+/��7�$w���5dt�����������
����rXƷ��)2��6w[/�a`K)k@Kܸ�<�u���8ǔaܞQt����Q�[t�����|��U�4Vy2�x"[�d�O�e%�-O��ţ���҄�������l� қ،nT���K��ӂ�i��F���(��� S&�V��|���L+�t��\�f�(k"u�X�� ᚗ��Mn3�0��^��@+Ǿ~��[s��� ����k%Ȥ�;���~=��<��M�H�h��|{��`Y�����&��P��h>�N��? b��6�h�D��6��6�jp��,Ӽ��,�c�x�4�1�z��O`��o'��L^�3k{K�M��X�2�ع}#���ıˁ�����<~B?�e��k�昝ҙ���:w�́5\Bve{_���
}� ��n��W����,i�s'a���G�l,7�LIlC�{��=T��S�쩸G�Г�	i:�&1R���I#�	 �hG�{��a�t���/�S	xAr��R���<z3�A1V*
l,�p��^�#�H��5�O�n�FI�;�U�
�
��5����V,J�ߩ,��>Fi'څ{�½����#J�����2$J9�~/;�۸g���;���>Q�C�~'��Λl�u�_��r$������Fn���=�ι�����Aq��Zљ�&9�>�\j5t�R�N݁��F�!	`�}�Â��y�n%/���q9/Q�߷U�R��5�X�
:U�BX�sjS���'0bW�%Kfg���Tq���9\�NR�����EkN�- � ]���2��|;��'�Wvr�]<]R˾��Kٽ��?c��=s�B���0��CD�h�+�M"W�g ����1���S3��N2���Bq�ξ��H�S%���`��vL�J��N�x���uٝFw��H���<�^�"2��5 ��y���sf?��5�F��YLY@fbh���z:�-Bn��ƨ��W��4��g��8{T�R�Wo@�<��|x�U`Ä�oM�[C�Q? �D���������cI��@b$��z��@(����W�v[8��ͽ�U5��2��E�+H��XEM� )��E��AF=.�	r��J�(�R���Ne��v��u�@����M�瞀j;�:}��'�lX��Mdb��1�Z�o�#/뉖�Dť7�������Uͨ��