��/  ��}c�G9�����~&�XY~ߒ�žV_*[6�y:���.�عfkG�JF��_�mv�UXJ2��r�Y��P�G�`=���<[Q�� `��$|\1�Z-���*��|�٪r�"Ŕ����	d��ܝ�3�d�P.-3졣jzW�2�25�@�^��<�J���6�����֕�%��!���3��B��b(�C.���3��R�wX����e%���r�JȐ�յ'���Pg�Ԟ�f�DV�	�}
�(�U4�����p"������b�`���a��3��G�&C�O����By��D�A����3���Y���_������8���w�}O+�BPt�]8WD��� �]�_f��*�(���,LP�0D��ʵ�ȳWsXڂ1�r�2��c�����d�Ѝ���#p޵s(��(pR�1�3�}Hа<ɒ��b���(w�e�DQb��~ӻ)��FP��G�uE�6}J_�p����VeV	ŷ�[�yKb�I���c@�S�[o� >�v7Z�>Ј�qm�\��A#�h_YD���W2�C�pq#)���c�u���,�:DT�}���T�����#�f
�f��=�b�@�Ԟ�L�p�8�;|j�	S^�d5�3������B+��Y��Va~��n$�Y�{�8e�u���/�TV�~�E��zߓ�lq寐��7��p��1E��]���9������O ��î/��a���dQV�ewɊ9�*�`��_�j���f��; (�wtW}s���hCBg��*�q����U���P�b1����zK��L���PX�/{)�6R�)5�ٮa�J%P.����=�.�ηwJ;H�?$�
'A�ԝm���R�T^A[���ɾ{�¦��|�҂g�F�+|�
Q|����J�H�*���}������,1���5��@r?�����w�t~�%����y�/����ه�(~@D(W���U�K��s�_Ea�j�����X<a��kg"���,�۠p�u�'D���	�)���u����"w����%S�'�A��.IZ=.a~��=��]�w���� ;Aɲ��y�?��h�
U'�B�����R�@��x���c�֢�SU� ��=��S�yI�G?���u{��ˆao-�Z�o�;��,	c��s�����-8�����&��OV�Q�}(|���f{��_��qx�z9D�L93>+�W��]�胪]��j|��Eф�\�XԩG�6Z��n�j޽t��vW�����aE�\��+y�U�(��@v���͐���a��;.��	������_09R, �۶�3`H2
sC�e���a�G9Ewc��?��V-v����OS�_8�8	&�ߴ����{�K	�l�\#

�р�-�����A�Pƶm��`����浉Xq[�YC2���@���N7o�z�&�PU�%��[n�r����t�^M�H��q�h��k��$�=H֔�#���ް���R��dӆ��:�ZL���ٶP)צ���%?�1�����iA�g�#���>�c+�°�'u䑩WM&X�N�K���N�ڝ5��ƻw/3���b+�M�ǆ��&vw�t|?�����d Ew�������7���4�X�N��(��v����Q�>bP��	1�6<m�a3ۥ�~9�-"џ�8\���w����`]��J���~��u���[hUΉ����H|騔������������a��������$\:��o�;�d@��U����O�G����6#�|�
&H���<}1�U�Lud�[��{��=	!ph+�}���,���+n���#Df�������Ѿ64��%Bt��@��L5�9kA���xP�1B�K��)�-�ɭ�@��Լ��9���
�p��5�9���e�"���@Ά�����iƵ�{�~U.�J�dJ93-̯u��Q�Qs���V���Q���b�'���ý��a��1b詾��}�V�G�%gߝ��e.Y��YY�xm2|2�]��6�>�E�+x��ٞ�5�G����5}��G�ڔ���>��=ƧJ�́�J��t�koZJ��� R�Q��-�M\�
�8AX�}	A��)�����h��M��_:�:h^#�̏3Y��j�!��;xC�eS�}�������>/��g��h��'������� ��?VЦ���z��5�8��&��n����D�4�0=Q2M��Ї��4��w�_|����b06���U_?�m ���Яt\�A��^%2'���½��[�(�P�Xł��Y��P�:"Eg�����5���{��Xkhp�����{jh�����o�l`kCg��m�`?Q�-5�8?��v'��H׆��4Ҡ�B�Z���ȍ+)6p+K�Qp��:�|}�ՔW��x��N%.&�I)���$MV�W�9�U�;
����0X݇;Ed�lݠ�^@k3��ְ���N��7J�k-_%���Y�����#�S�pWy^����w`�:��b�Hf���`�z_��^
ﵛ���G���B��n��+�?2M(������=����80ͽ�3&�^Ҏ�#�u��֯�0�M�9�p�Z5��
e�Z�q��2R�j���aiwۧ8gR�	=��f=��I�'V_�"�u�W��Wy��x{Wg5Tʪ�pv'�x��|�������U�ivj�vDW�M�8��=y��2�g���e �"�-�PLS���3�W���CJ����V.���\�����8�W
����_�UO�Y�oח��'(�����\wJ'�@�{׵IN�N5�N��r�ӏl�b��`���铭h�&��0	�#%+���ϋ�b��jnA����y��|���ǒ1�י�'��^�����a:��I� FT>D��k9�Y5����#Ce�kc�ʈ�!>l[6�l�@�l3�,�E$!1c+a\Ux�Z���ǚB���V՞��U<'�qa�M��?~������7�Xh�X\r�l����������)�������-�\]��x�'��d�?u	
ύ�����B�(�^����M�K�O1���a
+F�y	N~�{��Vq���E��51���6���3�L}���}槍m����O�ԞF@=�n*U	�L��9�XA/��������zC!��5`M6&�y��~*���>L3��B����<�+�����~aB��G�@ie���UM���Ы������ъ��#�K"�1��9$9�?n�?�K�����H~��Z?����PCǥ��y���U�6k��m/c}����7]��iin�GV���Nੁ�\W�����4�`�2o�Oc�I��܇�~@����8�4�Q0� ��z�p>�v.��i�E1(Cϴ|�)[����|ʖ/� ��z1w�g��g�F8JM����hҒ�2+����e�ӾF\f$�Lur�\��5L<|�>xM����C��A9B!f|���נ/<���4'?��:A��\<?>6 K��I�y�3�w�kOkp{;��%�o���S�(�u�F�nձ�C#-}O��`&�H��<�h��������ؔkவ!�S� +��`�m7�/�����4�u�U���L.�},#�\��\�!�6���÷�����*�mXMTd����I��_,\�S6�0@�~68���r�c����M>���t��8~���RB��6�i��E�X������D,� f>���D�Jmb]7=]SG���/���g3W�ޮEP���˻ȅ��Q���*g�\�ݤ�8ɓ����&�hl��/��=����`.�t#�r��~8L�FZ�Z�S�������jݜ�@iW��,�G�����"�S��7�EY_p �p�ůY�΅�,kK}U3���{]&�1Έ̕�	��+���KR��.��H�W�k�,^�I�6��o�=�� *�!Q�Ćؑt�X����[+�J�3U�e�=�Ei�%�E�ia�|bJ�!L|p؄/�.�q*΂���u7���`�� �imw��uϜ���I��:u
Z�$�<��ْC����nn(Y�#2O�O����!��bؖ�i�롻�j̉'|�X&ͯ�r���Lެ��� B)��4b�`��r]��0�.�H��ɌV%]�`�����)aO�cB�F(x؂ߧ?:侽�xxL�'�T� �,S>t5.@��,Rl�X����>��,���^�QKڤW������+�C�3ɘ�������·������Ϧ��w�Z�BX<�H'�6���.���I퓬���~W��%~�����Ƽ�f0K`��~:����Y6��Վ��-P\ q�6�	�^3�i>�߅��2*�E����J��i�b$��#\����7	 2À~}�0��!ng:�Qd�t��L??6^�7* �d�"�9M��@�c��u�4uO�0k�o��;��n���`/��Er؀�f����ڭ?�2�w{�-S�FG�7"#�YY�V������;�Xg�Ǽ8��V�y���\BwI;�l���9���Z.3�����z�
�y=YA�F�$,jPTRf�q�� G��^��u�V�����;�6K���
�(���sb����􏞑G�b:Z��B���t� 	9�ޗ%�gp�^7��S*H�c�	�N$).�鴄�i���+�W�_0�2����U���rw%tD��/Y���% �S�t�p3�#D�x�dIf�)��0I\q��
Αҳ��@�R�OE���-�� �cw�#�8��"~�\u4���!T
��)*���l���:F_��S���q23�c!��f�ւ�W�QGJU[�_2�i�_���H���d��W�K��^fl���3��>$�7Z��{E�<`�Ek��4S���4�%�����n
p�4�+Ş����l�a�2q6W��r��kB	;/�c��)`�O�{�-�s���ē]���ʼ��ss9Y6ߠ�����dkyq�d�����Z���Fv�"я�5�U�VyЮ��I?E�Ʈ��3We�k8i�$@}��m��v�x'�GqU@B�D�ڧ^ڝ�B~�K_��t�˦�G��cĸ�ЀW�rc�&����º�ٽ>���%x%D:��x_[�3/��Ř�U�K�k.��S�F��
e��Y�mԢﺮ�αJ.���8��Ю�"� ��$�+G� E�#r3t˕�%R��A��"�Z�8�b�6w�^���������X�K�� ƿG���yN(��̻O�0l��֌N�]'��Aȇ�����xf�������#�����W�(���P�t5,�$*fc�����cNF�\>���G�G�q��m���1.�P'�|{y���ʜ3���"ȃ����Xg���Z<jg#?�m7y���'�kbC�h]@Cv�x��ǚ�|�!�h�E6[�_�i���.T�>� ��7���U�Z^�e�A�! _
�p%�^3'�^�o���	���)ˁ��
ɼvY���@�ǎ�B=3s ~%q��0����oZp��/�w����1�h��qk�H�؎��;�"U����t���E9�T�>��&�o�-Ǣ���!�<��}�/��\�i���*���U�@W�@澩2h��΂w{h��)��-.���uL��Mn*^�^W~[�,2&ԧl+(��h?��`A����nL������(cIoJ�$��1#�\q4�Gz������&X/�P�̛9���US37 (@j�{sSX'�l�ү��N���rd�q������Z����ivI���Hb?.��7��U���������Q����0$�@���?�t�T���1����C6l�:z��
d���,o��ʙ�N~5�4�^wxo	x���ruS�W�z�_���y�ށ'��3��C��r�UFng3�a�X"�|�e����`yOΓP�U�r�X[��?�nS6{8t������?n��%�p��Ƿ��XqF��Sf>����VD�2�y'|�|n�ې�;�%�
�v��Z;#!K�_��5W�O^�KˬiL;���U�ԕ���q�5���g���()��dڃ�0aʋuتY��6u���Jh�y���ob��fh���(������꟡�]����$P�;�^�Y�N�����VU�Hg�G�u�������v�o��,�x��L�����艐�㇇3�:����{��)�ഖ�+��\0\�g�d��f�����75vb}oH�� (�7j�;���s��V!C�	���Nc'�zؙ�خ��l"�c�x�G`���\s��1��&�e�$^�����+A,	z��$���X�n�l5����|&u�Pj��͙�F�����s�A�;��V�ŋֹ-�dU�!\���11�ޕн�$��q�3{�4)�����v��d��\�3���u�Ԋ�؋`���XH	]mf�7�с���s����!�=]������C�k�S�^[��)ןd�%��@���W��}2ѥ�!+L	��v��\��!�״�QM�R�����_g���Z�U����V���ʝ��d�MJ��OGd\z!�ۻS�7�X�+�(�h�L��u(���R��B���m��2��
��{eV��T�&�k��T����'�	�DE��*��Gn.��w���m����8���K �~'p��P�I��S����5��n?\�o��`��U�UTQ�w����9���F&M��M������Ȭ�����@�IhfU'���HLvTSW6�u�kf暅0e!ϳ�M�k�m�Q�ȗ�[�/�lj�e�> Q=�Pr�-�϶�g�!�>{_�7 K���P��t���֖�.��|D�h��N?���cf��i��(T�s
��wY����׉c�Q�Ğ��S�aڝ�3@�]�� m��Ɓ��6�9.VT~0Gوg���u_͇���oq��?`���ăދ�����M��5٫�G--���e�k�v
g&�QV�J`�ЌЙ?G�g�]��Pl�X-����o��<�ԋ!�}�m�
��O��䥬pc�MYX���NY?��3dt���!Ip5X����:7ЇE(��wo���T&BSe��^��y��I�1�0���޸���-����{��\ZiGy$��%���-�F�����ʤ0Y�����2� �Z��|ã*��\���,ؔQ�XSx��@1��N��p@���f}�O��>�����a���zۚ�/�
3U,���X�C�3��9���SY�31q�D��xT��K�<B;񻁢C�6�b�&溒O��6�\l`i�96��M6�laU��2�7����U2{l������5>J_ɒ�8[���X�̨Ĵ����a)"]��:�Bm	�9<`���b�R g �����Q��z�b��=�@����B�4���i�p�p��晿��hb.�݄K�j����Z���9��U����+d�,�re�	�0�����&+���Q�^�ju�[��EE�MC!ʚ]�]���H��&��]��#`� =ͤ	��.�����k\���P^f�݉>�j��|���Q�;�̵������.�����B�h�i��^��M+���O��Y��
Ҹ&�/���C��g��y}P� ���0�,X������$5U�>�_��Q���J��;�v�~ό"٢���+��#�������-�^(�cT-�nq>x�u1�s�$�ZhFw���eQ�	sz�rN(�.��y2�4,{{C�D����m��]�LΦE��X� J�K�L	y����<�0o9�(ʶ�7�}Q@T($�mr�2�j'W�8ޡODK�ha��MG�d����
]޸_��GmO����ߩ�1���F:+�6��R������e����3*��<d����j�-ubZ�����"z��)<@�h㞛9T�LSt{�z���#8�_5�d��K�i�,��OPi<@�����㋅��0dB)Xsp0����k'h��(��P�g��7���ڴ�]�@Y���\����p��$L�H�	r���8��)Zع�1z6S^��$:�_�r�SŌ�N|)���wN�o&�56���1v�4�������U���k��زK�H���)��	"�#xI�z5�tgŪ��E�\G�Me��PX����o�ɱo��_) ^�H/��| �.[�Cv�+�L�,�x�����C���Z@2%髯��������q\�r�7�j�&���օ��>�R1T�v/Ί�]��qV�	#~1�SE�3N&�@9�鿘A[F�T�af{D����ؼ~�,��Y �	�ή�5L�w����Vz���R��ܨ�U�^Fs����7�z���᜞�C����R7-���D�t��F��S�~������܌��P0�W3|
ۡ���$3D���v��^�t����#�z!Iu�\$Z[�7�XJ�t��n��� H��ic^�GwZ���I��i|�g���nT$ږ��e/*�zٸLиn�LZ]+^u��a�N<�=Ȑ� �*0����$=/�0�)X拫��t	"y�����H4-ڇ��.�{h��V��*m�h��և�{����}э�a?��g�E{���J �&�!�����f	(3��">𓙫xؿ�a�$!�Y���:p�O�p\�N0����0wT{A��o�pF#��ZAO�g�X��+�pҜs{�1�7���o�E��M$�c��E�R{M�߭Vv�f�0aG?���z��>��ĸ(dE�� ���־}2J�hf�k�T�Uv���4x[�v�y$d;�}�-0'�I� ����Ƞb���M��arq�R ��)|�ɏ���ٓ���e"{��]]�H�� L���7�gb	\��oD�i
�`�-�=mO�(I�PUA�h�-�0I�! �[?z?OK�Ku>yF�_7�a4�q��@a�&O���9�M~�5d�j��P�єoy�.l$���k��#h��_lt�4�3�<|����JS7J|��\ψ�E�j0��XB�l���*b�M�D��+��
o��bp�؊��NS�Q �(��bE�d�[�
�Q��8�k�x��)�݅�,!W�8-�,��K�2�ʛЦ�S�R&(3~E�ǯ��$��<����t�@m�9���d�>�,_�%BG�,0�N
2���"�.t��baQ�]�3��+�*z�)��E�u�K��\#�'
��X���upl���=�����8�p������7�+�<��D��1&QIT
}��k�j�ek�'gl��~�p�0R��"�˪~`�
��B�+�''6H�Э_�ψ;����r*C��F��j9����!?X�Ƹ�y��L�E�H��<*��t4�|��Zs�u�)������Y8�^��s�9v��p!׳
3+�d�&�ح�DcR������y��"g�Ěݱ�n��8�6�Y��E\�q�e�^\�(�VD[�ݣ�(��zXg0jᤆ���4�)B2u6
�V��m��j��x�����?@���C��}��}_�E71 �Ȯ1��=�.�!�c��������)h��rG��Ӂ�I�05�*lUc����:�4u��ώ�x�����>A�P�d8Nq[@W1������"��A�ڦD��NćGK��إ4Bt��Pa���
y���rB�D�u]�=^��k�"�6gOyV�MN������8w�q�[���� ���Gu����_�TMai���AFkQ�j��6�����;`�ш�d-=ˑu���Q#cY�MSjl� �O!��^��ť����_
���3��H&H���F����Q�D��T���Y�C{Np)������� vXh��}��rS+�4�����ǞU�L�S��dCBQύf!��zƞ�fܝ{ץ<"�{�3}��{e��Q<�̨�Un]+c��#6�\���J�+Ary��k���FgU;xQ�
K�l�ekԫ�.���;s*-��xaJʉ�:��~�u�P�t �4�\A�H�*�rmL ���t����xc�W&��Ձ c�n쓟L"XvM�n����N�aGD��F��ۤ����U�9:٤��H@Iˑܳa�H̗c�K���h+� yL,���Ď�۴W}3��}MMsf7�x�03}ߧ�@e�iVT��8��lQXr�^L�3ǫ�> /=����M��[�P%���� ��մ�����4�0 ��� >�D�iA�#�Gؕ���пӡ�������TIo#�4|O��{;��϶�fG����=}���p�����|�����SN�H��՚�~QF���+��ۇݹ��NC��y�QGfu5ʇ��1n�i_}��鹧� ���6C�����P���X�w�CaN��8�j�x�V�o`�C���i�!J��klޮ|�������1;s�#�%������vC�2a�\`萸��:3�+[�x���U-Q�~� �c
G� V�>�^��?a�\�k�ѫ�+Ǳ;g7�~�h�����ޱu1�?P~�$��{���Y��E���r�".��i �D.��	�t��O�f�(��V��)3���ǈ�Vi���p�(�<�k#���-�Ҧ�a�U��Z�?)_Eā��a2�j�شg�����4� [�@0O��E��}5U4 *��آ��G��TK	�Q��d��O�#�51��;��[x0�7���	����7�Z̴Z�z�5>���VX���[=vK�ٯD��DU��Ñ������ݦ�Vf�v��}kf���p�z�	x؆�U�lӸ���*\��^ٝ�Y�0�6�F�1��~v���Kp���Raɯرe3}@uj$�l��G�X�*�DUn$O��~X�"�c�uZ~���|�l+S��-xW�뉤���T*�"���p8�h�Ⱥf�(F��g�Ȥ���"�0�B]bs<�\�L3���/���C5L][�k��G��ϓ���B��j��4y�<9\/�	.ձFd�2�<w^��G\=��ãV�\lT��H�q����Iu.�6�Ԯ��J#U�y P9[�\B�x\�X��J���x"�Y]��ն�:oy�4�֦x���w�͈ժ)� lG[���n����)�N22��v6K�@VS�>y�k�����qY����o��q���v�q'�R�2i����M�l3W5Ȇ ��_x,���H���T�shR-^�h����1����]	�)30z�t<���'�<~b���2�Ki\�k\Tv���9tES�����
=�`��Q*��A��2<܊R�Ol]�<��t�R�a��X������O��̾����@�3x�)]sya�+�{,�tW��9/��$�rX��i"�({�F6���/fK�pʄ?)8`���n��V�^��.�(�m�yc��N����4$���ԯ�M4�۲�Ƃ���i|RCT�@+�^Q�mPn�j{�p�q�=��_h�:A*Ϧ��(]
	"�)�#�c��Krq�.�� `a���=K��p�=`��.݂2�xif9�M����E��֠��:cP7n]t���s9�ł�j���5� � e� �W�u��gө��:�̟J�dz��Gs4-��������P��6f���h���������E�2;6��C\��K�]����f�ރ��W?^�㧅8m/yS$mC8��|把�����؞��|��	�r������]xSȸ;r,O�L�@���G�O��k�"6wm�����k���ߓ�kpy6�r`@�jZ/ج�w\��G��Evs�⬝�����tYm/��K���i8I˂��u��gg{0��-hT��M2���ܪ���4�v�(z���,�{���8��K>��	4V��a�(�IJ��r$
T����t��B��|%���+������ڽ��:7M�F���5��|2��g��16h:x`(hs��'�w������j���ɸ[b�u�F8������u����M~(�L� ����}��D�d�Ʀ�H�Wo(�<��W��?��9f�jsWS�3pW�V 1��70���RJ�T�H���#<�������<�v|�&���ڙ����6�0�#���㞄g&e����.�P��"��M�s��|���U�x��a��e%�U�큡t_�����=��rw}���(��u�z�9�mh��^���)�d7����
2���t�Z��L�E{�h��ֆ�X�"F�E#� ��/b��*�^�f��YÀC�������
�����`㤜�F�;~�߱������	9�lN��Gz ni�z�iKr�֦o��5i�����@�C�R؇�j��V9$@����������?퀦1�op��~�*i�D�� �$��rk�v�Vd�=�
�����stY�u�?\��Q�h������0z�i�_�wsENF��f����p�ǽVVC��&�y5#�:��h��F��ф$�xG�w�	��W
�,O��u�,y��#�����iF�k�٥��P��B0��?V~�_A��X�f T�Ґ��SHe��wzd���M����|y�ѵu�N`�In��W{��޼�}N��Ueqۡ��2����b���ۥ�����:._6���u�-�uT7=%�{�i'{N�u�o٬�i�9�ϔ��r"q6��7�?�t�����8~�Tè�m�<`�ސ���ZP�E2龥��M��X���<r�q��{E���QJ�&bcV�T4�%5���+q��N�Ie�%�D��I�8�t;����Qp�~���TOƛ��oU���<E�qy��~>��d�I����Q��9�	���	J;�B�@�6���2;���09!|����t0��T�(�v��r��Tg�9�F�IM�q�3ݰ�<z`��Q��|���$�M�1/�Fq�Gz3�D�u��U�K�$ldL:�ݜ��z�hvڜ�&� ϴ�G�,x�܌���*K)�tc��^XP���?��h�lk�C�����B���Z�o��ZV�]�Y�4hq���7;��,�p��r˚S;����+H]c*0�ʪ6l�L5���{X>�<F�f]�`���$@X�n�+OE{����a1��;;2ʏ��$kl����`yǸ)��q�v�vݛ�z�~/�e_P;��W�H�����j�w��4�p~�8�O
�<r`�'5
ؚ��;�Z���R���U���BZߚ��H� ��t�������;�T�k��¨�RiB[����Q � �#J3󝦝m��S��&e�{���а`xU
o0��2[��p/W��s�$w&[�� p12`'�q�&7y�2�Wt!{ �V7��o�o�cԬ�G�Ci%��?"V(�,��S5�3zF2�dr1�>_��.��Xe��iK�a�3���S�ƣܳ�E�n�hT��f���l#>����!�����d�ƶ
�[#�,.+^�J���p3��碑}s[h��R5�j�ΉW�M[��`AW���Mp����0(ێ!�=�*�s�r?� �M O��Wg]<��M]a�V֘u��-a��̒���~�N�{(���O�E���}і���kC���ۚ@�YO%$P�g�tf���E��Vq���>U4���ExZ����6��k_�N,FP�;ϒ#H��(_�K��U��!^��,��ݻg0x)��C>	a�h��°\N~��@y���;�=�f�Oӛӌ���.I
�މ f�En	4vΗb'߸=��h��(ٞv�W7!�+l�䚎(���{o��'fF���xKJ�IE�;�ĨU���4a'�! �d)��0۫u(�*�PG�Д�*H��p�R��G����7M����h#���@��t����j���N��0�jj�SN�Ȗe���1�M��hIG�>	���EV1:o�����Aw��s�3ue�ak$T��鱃&}o��n���+/�)#�%����͆>�!�d�^�$"9{P�XC���
��׃Cbt�+8�2�Vܸ��-3�T�V�σ�=-M��o�+e�b���v?OtD�j=2�\�1�-
�6��4_����u(ȿ��P��qmD�kN�{�u�e�؀��"?�8W�Y����l2�h�si�8��غ:�2�=ѓ����5R݊3I{blϐ|f(�5�[�D��8��Ĳ5r,�[�<V�4#j�`���p���w:�WlKA�u=��,`C	n����kD��,����]�$A[�x�_�4��Vv����"zG�P ��	'���ź.e��.�~0����Y輺2�w���﬛[�ø�D!y)ϼ��n(���l8�E�i`˸��r��P����&���g�3��|���}�@ˡ��IV-S7f���a�_f+Pn��<Z�$��i�o��ŦϦߟT6��^�*��7#�����܁pV�{�����a HY�����C����V��������ҹ�T^��5_Ń���S�#�a�۴ϕ )��z���:�L]s���'rA/����z�m��Z��q[���j�S!�_&���n���0&��ڎ�9�a�x����&� �e�����������8�9=pQW�-��$���ɨ�e�D��j�~�%]U�bd,��8J�C�Bqp���qvFG����/�Pv���Q�SE+��$��I�ER�*�����ۺ��Ѭ��w������	���9~�m=�'��*��+aˤ��&�pd��C�)�����_WV�b���mſ��ﲻ��,>�o��Za�s�R"����	ЙE��v��Vǳ�k���Ƞ ��U����v&�^OAd��h�ÌR���2�圼�s��w�8�_�x���TK�)9���YOb���__!PGRT�.<.��Iڮ���.�Sd{�:T�fq��>��Eh5S`@��0hv_ӟ�K��a�~;�f��^�qa�kܡkd�_�r�"B��T�v�p���P��2��z �Ƿ��a�e����aFJƮ��B�2�d[�]&[��jV�+kt�e�B�l��$�n]�z�TLd�ξ%�t�F'�?ބΊ���{���(�5Mi�Er�7Qai�L��,/��
�Ì��\wze��PGmx�0E݂��)w�� ��w)?��΀���Hkl����Y�bG�?��g�o�[�p�ն��SVTz�7i%�}xh�|G|��jgM��= �"0 M�?���5�ԛ��ך������|��'�g���j����蜲q[:��[@[/2��Dj�L��b$�{�7K��5.'�08�gq7��J#�R�G8�� ���xILگ���ȤV$�c�6��"��I�K�n��^�D۾�`���O����`�|\�Uc�n���@=��1���:
sB�*�ًۗg�+�_���i�a��=�Z��h�ȗ`�E��W�[�AP�\�0�~�Q�ں�µ��<0��U/�>W�\*�*���SM{�SA���U�c.�`�[mb���l姢+_D�U������.��<�\o��8ޓ��<V)���_]�1[#�%�u���H�(�2�@g����_ ���(�0(������H�"�]/!����!ܡ��9��6L��̛�!��)���&��(�6�:����SXA�������p��y����Jk��Կ�8ʘ�l.��t���eY�+��]2�%�@"j#`nv�HQ6���@\˒dH�LN'� ���"�*��ڍ?�7YZP=ˬ�1�8u9�����.���(���� �*[�j����
y�"꜆c���%6��"J���7�u���Jx��3�E��x$԰�/f�b��K�ti_Dme}eE(�~q��>�LA�/�{˨����PMr��ا6�ꉹX"���U_�o�[�/s)i�e-��x�~Q�H~K��G��f����7t��Ĺ�ˆ�l���(�G L^O#A����C�-T�)Ea��r�����R�.��N�__-UiO��{^���C�~`������қ�A���[�������$?���ޙ=�ji����k�^�ueF��i՝ ���� �u2��gO�r�����sz�[gm�H�8� ��i���K(S��X�TBh�P�i�q�1����?�͏�2l�ouD�Q����߶y�t Oi6�s9H�}R@-���n��f�9�]���^b�Ή��t=�/@�a)=�u,T̰*6�ޙ)uz۵��r@��y�|]L6��������<4K!�/:��u�DU�G�ˎ��7�$����� �dVaG=���'�7�z���EF��e�|sڭp����񊳃���C-���tɤ1�L��Ɛ}���FH�%'kG����qհ�$^����q�?�)m�XcQC���(��w,��v�8�ths���YzӰ"žD\설�Q��'â~�&��t-ĔRr�����E,c�80G�#��z�j
Ӭ*Z*�ժ�'��7��4��B�"��l�p��r���Fl�����j|u��=Ij�yI��ǳy^2����GP��kA�{ժ׊�ƻ�ʼ���,���k�>�et��{qF�%05\@Az7����K��T+ڦ�Z�o��̢b��\���b���T��T+��%���徆pTFD�-ʬ��_x&����`[��2��S���X �\B5����h�K�T�M��W��%����K�JBy"��~�4��D���l.������@]��Z�c�0JuK��kQ�u!Ϫ� ϳy�P�(�'�D���GQ���3��'0v���CS���+tFݕ� �K8�Ta���Gr�����=+:�;��@_�S<�I�{�&|��~�U<�}�8b,��X��#���t�@�3#in�6S[��dZ����6�i�x�"6���Z��O8�����#<�bqvW�Dr��8�1����.�lDh��V�dzF����d���pt͎>��]���$�M9rd`���*�Ը�MS��	���G��99İ��ڬ�>���g9
{:+��5��A_����Mh*����c��d�JG�y��mZ3����4���2�A�=��B�h>�V�S�T���?"�7���k�?ey[D���#��=��D��_��}����/9v)�?5��B4/�u*�49���@ɶ�����=$A��t�a��D�#�����]z�t0ۋO�����$�F5Q��_o+pL	�g��!�� ˣ���F���x�74�˾��Tme�u�B{��˫�x+12@�.;�� *n������O�`�џ;U�"���#�%�:��F��# m��%����i�ĐsRɗP]�<��9[r	�h�-$��+~W��D��f\w%KJcf$a������O�pB@��R"�]��(|�7�ՖnO�o�Ԛ_�&�؀�Ki$L��n��EB]�9����v��~���8��z�d��j�p�a:_ �kJ���g+o�S�\�hYŽ���R���bu_w2B��)�6Q��
s�h��]�2���Y<wHҦB��Zb�)W&H(O�w�? �S��?��cl��\����[;�>
Y8X$P�q�Kv'�л%�<����AfXn�W�Au�<����,��?Rm� �Bc��}�,h�y����bE�{�z�*��y
)�D,7?�P��a��B0�V{U� ��6Q� &�B��Ϛv+�Q%���|�G%���9���u7�E��-E���iS���mV<Ϗ�*Ϩ���$Һ��FF����fr]>��dI�����ՐksQgV�� a���YFj�y���<Rm=�w��!^�E��9Ξ@��OҐ�:�c̘d���Q-��p�ߋ����Ǵ�v�}C��x)ȴ.d��.�B��)	���i;�G�Q�qns�bMv�8·�6J��SV���\�9���I� ��B
[u�|�b>:m���*�Xd��k�<���������F���r����9�_eZf�"+�+���$��;E�3Q�;��}�,Nnjj�[x\'���u��o�pgӡR;ʓ%~�����OIZR�h,��w�6��r	�W���x���Wc����'���%Y�n6߶	[`*�*C��h�N�mR(��A%�� [�Ν5�px�:�ڿ�|�~�9��:��a��Ȯ*����=��޿�w~��t�9�\�^��|i=f[�l���(̠	�l� {�Q�S)����Q���D��*
b�.
6�L_��|���T�W�4�r�Hn���ZN����:�<�Z�2l�n���z�lN�@�=�"	ذ�)ci���POf�T҆�Q�zI�>Q9�}�^�NG�'#�ƲhR%���K)�n+�TڭW��[��v��3AS�X)��Ё�O	7b�" ���&��+R���0�H��I~OX7��K��r���&>ch������2�Y!7�����涾�6`[�j�B��9t�;�%4�KU�.Y�>�͑M��[�_怠2� �:�$Z�v��&D��5��H�P�|P�Ov����������	������$�s�N�>���x��7�N���
2{_��}�M%�;�4��1������I+>���q�9�2�݄`��Q��Y�=Ȍ��9ܷ#�4!�܌G#�!b��'��!��}_��4�iP:�
q
f��i?�Y1Kk�^�haʾm6��C���yRy<�V�1��I�=��C������crw�b����G^�X�\��]���|���e7�K�HU�,8kZ�6t��1��׸e�?,3em���Wh��u�^��5�7���)67<]�L��ء!^z�\I�{����@zZ�N�|��:T=�-�k�f���F�W�|�Jf2����&�O��U
�h�p��YH�-����F������Y�n��x�)2te
���Y��RQnuqݬKm~�~�	)�~`R���G�~���!ժ/,p�?��(�B���Z��ct�u�E��l�	J�n����ـ�v���"G�����|��vmh�6��p#b���4�
��\�S|��ٗw����D�I��>l���nL��r��u%E�&�fk�&W "�<���Z��/�v���4�.�%���+�,�Q����D�$��:u��t!J����[E?J��/i�5�#G�υ�J�4������=K�����v�
+�T�I�8�y�R�����(�~C>��D$�@Q�n4�_#�q�������3�a� �������?����~�H����^����w��h��p�~Y/�vx|.��a�2k4Ʊ�S:��Z��C�$NtUJ�yҙ�';Jjؿu��Ԯ��Ը?��a�5�)Bf�;{SQ��:�}���(˵���[
���vA���4����E�6��aՒ�T�B\�����ZV�>8�\ΈUIt�ѱD���S�p����z�ش;	8B'�]g�"b��@yz��mY��	Jp����!�J�%�����H��~��G�]O:�mE�/��f�	lM�_I���Z��qs+�MQ�O�Rm@&�'���R-cXu}BA�}�^�����SM�ik� ]�Ѹ`��q�8Ϳ�be�@�-�~Z�Ֆ���9T�|�tT,�$�Pu��~����Mn�7+���9:���� \j�����F����p_� ���h
��l��+�b���lm�*��r-���U��ޭU�>ˡuN�Rl*&�b4��Z � ���fʅ&�Z���r��Fl�e�:���tDxc:E�.�� OZz,�`5��5�����ӻ�e��e��e�3W�`�L�^uCŤd\�V��D��-��o�q�,v���:��u�����&<ɹ���
��t�i�_FX��������F��9��f������o *�I�	h�<�#K���oa'fb��g�VA�I.�:	u^���_�����tA�?��⦅�P��@"��tu�UIe�}W���n@���j�@�;)�c����94��wZZ~?��'�غ���9��2�e	S�է��y$[ί�E�Rw�a��~���5�*b(�y��szgv��߉ɷAc&Hf��h��<�[�� BIY�4�L��RGNK���x� E2���d[�������`� �P��y]?8f$v��2�$�Kݎ����Sˤ���t"|~��@�����]�Bw��iHL15����m��5������ƭC�īh"�]l���ц�N��w@t�[Bt7pYeC ��7E�D9�1�>��A	T6��Y�l��1��W�����N�XV�t�tiWA�Y��f���a�c�B��]�aщ:�����_�A��-'ڳ���&�SL���!�%<���-HZK`�W�Ɇ�w�d�5����>P��L9�����g��YA���f� u9:V�!�����r
&�cי�I��{&SF����䗶2�d3y/k��Rl���}�&��f�(l������Hb�ȡQ�/�f�
�3 �`�U���m�V
K6��s�ai�:�D�TBm�����'����Sq��]��rC�'�dHi�A�Df�Լ8!���2��-�������d�h�BS"SR�O�6�-��T1m!��ґQ�������,��z��X<<&5U9 O#Xjh�e%����z<U���:R����l.'�Oz�p�"��[%�������	�o�)!�b������!��������X*��ݏ�%�(Nc��<�$0�n�/��O��w�*FW�q�8�����\t��%I�ݍu.����U�	&�B��Uʣ�j���u�o9*/(䙹�)Ξ^�Q.��c�x/ǈWF�d�VV��
w������Ȼ�l�����"�`]���4��$����,&�)�G�0.C#�ſ��q� /~�Έ>TZic>-�
�H~.�S�+��8�-��= �o��L�S ��Ñ���lX���� c,������Q�E1\#�Xk�����)e2/<h�UBX����"����IK�i_�� j����Z!�U˪V(z*~uC��a�����Y��F�}\�G,�2i�c3�Q�H~�l��M���V�c��=X#SR�.9�����L�k���0�Ht�ត��h/� �M[ҥ��ЬJ��;��Ճ}c�ܛ
��lE��:YI��<�$(�N��S�,��%���끛H�g��y޺#YJ-?��ۑ?�k��ヹd�N��͆��R~K����:�Ì�2cws�)=��%(���&��Û����wi�c�,F���i��ڤ|�g��wx~*5��#��qY��w1;L!&�J��f#�c#Nm�#�f� `�m�R��?��'���q�U4_V��,|č�e�� �e���� ���L�'�>�����r���i��x����pQ���6��@}�K_�f7���jkmJ6�g�'t7�
�*�T}N���u�-����O�s�j�ӤA,�!�Tg�u3B<ew���q�3���!�G��h��)��ʂ��˚Cl^������mt�e�	z8�Ī��^1�
<���\9�s�2���W����_K�ٞx�*c�Qv�Cp�-[F�ØoYԇ�M)��s���fBjQT�p�.��.�>��3�i�u�M�����F�EN�Y=\�ܨ����]S$��﫜�}ҷ�W�(9�}C:���nu�>-����cٓAA�>[6%P�K�y�$M��z)v簥�p��9��<y�0�X&b$��;���(ג�S��E(��^�������|�U_�n~T�����4# ��bLQoV ��b�M��q���B�վS+��*Z�}}?����]��<S��9D+A]����^�n�8��X�{fzp�-�'3��oWZz�B�`�}��I[��0�p��g-�����t=�bp�`T�U�f]`_L�\ؗ�i�r�nX�)�_"R�]��ҽ�c�cE���bI*"�`-Y�|��A����/�
t!⁘56�π�\5>���IFE�F�E��|`B����n8�s���$lK�i�}I��']G�{��ׯ��Djp�O,��"
�A��"�y�L�kM�s��/��z����<⼬��'q�1��c�r���&5e�f*��AH��)���Y��������!(Q�ʞ�2,`A�u�m�X������9��@��D�����e�ḌA���8gD	|���>mT�	��W�HC0��?_=��7�w�1�n�Q��֟l�Y�w<�������4@w���}����Ÿ۰pm�)D�N�%/0�T���,��6:�(���-A��(��8�`������꘳*���!��͂��eq6`o�}�s�V.����5���)�~��w��t�!9�lѝN��f�ʲ�(��y��8n�a�z�2�-PS��x�ѯ�U9:҇,�R�(vƝ�F��C���a5��@�c
�aD<6��"�k+|��83p7�9���z�����ڎpl]ȑ��@[T�O�P�ȻSOkL[�m/N�Q{��"�߃F*��!?	�
!�{MP�b�yq��``f��r9�ۡv5�<�����o"��D�dG�R��c�߫��9�v��Z`����r~R�(7���5���רKo��O4YɲrOD��&��x�b|X�s��na&�ކ����6X�^G*�c0K��60���J�!B�"�6L֡�7f
�iO�Y�hA�*��R�;���@����>l�#����=F��Ӵt���LlC��|�BF�ЮUn
�
l�93_�1WT r�0��V��U�8ʹ�´��|��p�;�s�p�+����=��u�B�*i�,�I+B��2���%��L'�X+��:������9`�>��˨����Z�ɐ���y�c/��+Ͱ�b��^c+�䥾��E��C�]C2����_�$����� ���>�h\�r��q��I�H�/=��	w���BL�t�>���,p�|�M��I����"���h��LE�AԈ4����Zx�Zq2HM�KL��1 "��%i������dQh�;J �z�
�d�*��`��K0̖iM��RRb�A��������y���F♘��S�d�{��#�ț
����?�v]^@q���_ %M�gٻ����Bl�;()Q�R���`)��j�C�D�(���Q���?Q�/.x��	�;Ϙ�Eܛt�}h��[�N짖7��q��o�K�r܂L����Er)RE�O٧k)� Daq���aD��FJk�8��);+[�p��'��3 �Zd'
�$歮�e����xa"n}J��cDY�8Cʕz����m׉NT��}�D��$a-i$^]m+i��|�s����G���G}�@�$�I���
m��k�HEp�ʆ�Kj ��A.����|3����~*x�+���I�A{�{�.2g�,�kLgȢ52ʝ�q6'pӷ�ns�cTT�;��ڲu#'��cބ֓d@��I�o���ҙGp��D�~E���]�����Q�y�xx�p����	C�K�)�����ɥN�&�!������Q-��&Uຬ�
���߽5�sp���*�P3/��
3�e8���8Je�i��������S�	�����(i逎���o�8'�=K��db��N�]x�#h��pT�ʄJv���e~�Ž�
�,�&��� g�@m�4��9\�6�r>�a������NX��jm'��+�+dDlT�)r���'��FA� /���錻��`∢�TF1�e�<�Y�k/}��
B6��gkɵ�m@E�f��-b�^/��y�~|t}<���[Alw�q�/��(�V!��m)��{�EXb�ڃ:�N��C�b8�v��
YG����d<��!B�.}j����y��&�:�!�A�йzy^Ӎ�.�irr��y��Ff\���m٦	�q�HnO������'&���:�rj��Z���� �Z�K
��/u�K�ؾ�GG6@�cϫ�O���0�Y�@D#ʴ �|3��3�\�H����o�Vx��l)T�U�}��)<�8�jMҙ�	�U��C���t�^�I�������ͧ���C��O�`�D����#�YJ渢Ð��G{�}�@`�p�>Е��L}�����=o�;Aq���T���Q��д��.9*�;V�<�̼V^����Y	�������|���3����YQm/>�)� ]T�|�yf!�`iry�h�F��
�Hzىk/�s��$M�q�>�����{H�jf(Uw���䇼�����CB+�+���7�z������H�Aj���:�f��Z�.<g�+��KRS�`���5ip-�s袇�Dպ�Tp��/�"ǻ��7z)q�$ �-TKUu�cD��v�^�U�~�.<A`K�H<�;g� J���T�=+Z�������.�<���;}�V9�48`X1�)��\���isQb! ��m#X|��m��v�[z���ߊ~���d�� #+~�;��p�֟�о5|�_��c@���W�5���=B��$zd�o���ʍ�=��H?_�P��,'>�ɢ�uώ�1���4d��,��������^��u��U��FeR*砾��{c$3��z��0�>�0�0OU �l�LFm����`�D����QK���$�1�
Rm�}�\�w$0B��6l4�9�|8N;���3��K]�����ú�	[��	Y\ٮ�ԑ�:G/��>�AI�{Ū�&	`ݮ�9��V��>�%��z�׏N��H��=�K��M:�R�a�6�c�K�?��K�K{��h��;l�]�M�����T���m�R�=ܫm��lov���U�h�nG�]/�Y3�+b�"M�u���e}F�|� �4����1�2*(l��|/XK׳����4B�q(��*�%#�漧n�^��O����7x�d ]�E��A|�4��w|�!��VQ�e"�[���������<�O�_ny���2��2��CiY�SH,r����q���������� iP��E�Ԓ����E&�c�:��:�: �ߴZ�n9�#[[+��L7�=��q��^�\��R���W�0��x��������V["���
�_9�ܖ/Xӱ�c��1W�#RW܋JaHNBb�7���*ʮQ�,��:-^I��p���O�IІ����5V�{Rl� /A��c�ET��wI e��{��Y�6.�(6O��b�t_^��e�x�G^��0�Kd��gI���T�U� c�n�g�j�����rI;���הϹ����)�~~ T�xV��[���̭,|��h�=�n�M��J?
S	�k>�^ 0uO��(]�~�O��kj�D��P/XjKe��װ)�:�qE�Eei����T��� *~%R�N�%X]�Av��'��n��dt	#��U,�~�R�+��?�:����0%�f1����8$N�;�Q�v�W<����~L�1�e�}m�@��B�_E��Z�w圇��㔴$~+��9o�{<��X�,	H���^��+�ۏ����,~Tt@bEB���K�Ao6�f��:�#|��d��5K?�^��%l���D�@�����T{��k$��qj r�a����gl��!Ǘݎ��k2��9(q�7@�0KҠ���{�<��z��N���b$�Qr{�xD_x<�[���:�%�����B�]�yf�3�Q-��OꍤѱFQ�s��x#+�}�m�P�\֜\�� ɽ!��k)Wp�}�ac�c�)��C�weV�r�]G�z���	��n4K���n�K4��V���|�=�Lo�,S_E�[�s��ֽV���,�W70�g�5� ��|�ߧ}���R���nR&�r���ۋ$����>_Fn���ִ|�?:�_�@������[d�bԺX�k$7����_'�:+�>K5Z�sTAI��8�?�Y��{tG��\��$����d���˫��C캔�������iS�FX�Zf3>�^���
�^��i(]��Āˊ�p������V��o:��E65��h���٢��r�����z�*Ɛ�e��t��y���*����H�Ɛ�ZC��@$�B����;�<WӃ��,�f����:�
R��Ӆ~�Q�ez���8��#�%2_6�o���!Ѽ��D`�7����L#�+������Fw��]���:�ˬ��9�	W"�(y�p�I�`���i�'i�̪]A�cQr��ŏ�w��E�)�Rl�m���⦬���'�������<+TF��9�oj7!f+٣�0��Ww���:n�� �Ŕ��P��n^�6�VaZ����\����Z�р�u��������-jĲ�(hN%T��je��OJz2۶�������[���@+��ؤ`���Ӽ|x�.Pf �����!��%ѳY�[�TY����Ѥ�ط(��{��Ϟ����",�K�U�н������<��%��MU������׮���u���sMK�t�=ox�݆�n�)[��$gC<�n��
Yp;����DDPͽ����q/T}UDT2[:n�M�2�����k
>D���'*�i3����K����d�� e��Fq����e�ߤ[�z5���/�I������|����bm�/+�ay^�wɕ�̕L���/�C�����T����}y�^�\����/��9�d��C�*|w#���'o���Iv����_���@��Ե���(*$P�lC§6%��Ra���*ˆ�ha[ЌI,�ՓC��8��A�P�V�hӹ
M�f�l�@��dw�c�gk�Le!J+:[U�G���kzT\���F�D�f��VP��q��h����^R��(�<�ya��S�h�9�_��'�4��6ڟ:���R�!��	IR$c�IM�"6�#�`<�=�ߒ���B�ᅂ�J�D)`!a���߷���f���9�y ���t.��[����sWX� /&H�r�8_�����G'`2�O�c��@�[Yw?�AYZ�"1e�Hq��%��c�tؗd�z�<o2d�u�2��25 ���ԃ�g�]M���ɏ���Z��2����g��k����X�����ў�;�ʕ
���_�kU��N3e7�yEH�X�\�� 46��$�F�_w�v�X��^x4rL��)_Yޡ`�9��6�"�$a�k�t���QBޛ+}���e����O�]69v̺���E�H�]6�_���K�]������'�_g��V��많�#����7���=:��?���l;��[h��U�8��-7�:4�1�JZC���e�F����������w������ϴK�V�6/�$��^��5�����P�g`d\ёP���ٛ��Y7��wgm����%���^�*�}��KZ��͡je�B�~-쏏���L��3ݿ!{��O����"}�R|HH��fr�`g(�l�#}�#\��Ӣ ��I���"#8�qM6�ƫ��fD�@͒"Z�|��H����N�C6hl���e�54���Hs��A�[��ɑ���j
E���%��`��^��JH�Fb2}FVK�������ń(��!mܢ�Qz�!���6B�ށ�hU����_��5����vsm7/�FY��,D���e����Ĺ���(�/çUC�c���ïJ�,�m�ÊKÀP�;����P�����$�����+C���Ȧ�C ����2YhJl*��G�6nU��K�)���[��"7��J@3���^��I�����
��P� C��Z]�q�'&��2���r��y�v�(Bl���2A\M��/+$��W�.�8��x@W���*v�
{%qp��c�>�N$Ex�p��P�mJ�-O%�j1i�=�{~K�"ò����U�|�eI5��'�#:g���Ƣ�*/k�ƻ,�_VO�i�<8��e4���aʒ��E���7�/N���E�</!'G��x���/c���̭���g��R�뢕 $���99�8^�*	��j��}0�$^!�
��� ͛L|�)F0ť<kA)��Qћ��JIU���:��U������k�:�< W�Uu҄�����͠x �m]q|J6���i�)���}t�v���X>�G���I�Þ]9i8��ݦ���=��6_�&�[�J��y���v�����P]W�>���kII<���	�p�<Do��	ď��Kr�/������G�1� P[NtE4���\�p�h���W���K�Yt�v����z�g[n�䳿������{�K�c�/1���8�C���pKoЉ���x�ēDϒ/�#�Z����K�������UXxVH�\�?�;�-�%�D��ɘ�*&Ɂ�2=7�sq���N5ep���Bn�����𑠹�a�k��b�ư������{!Nʊ)a�$ P�(�g�ka�<gU׳>G\��<l�~��V�|��99���ꮫZ�!������x�)���ԙ����5R��f�HV���N��F�I��fAKbb��sU��R��>�-č�_
EuH@�
�yRͺ⤚&;��ϓ�&K�+���t�}��y��鬪 ��֜�K�a���=�\��鸅u�������EW��InL;�h�%�(��k� N�ޏ�BO�%��@9s�Tʈ�̓����n�{p���" ���Z��9#��)��]~����߭�z�&�n3��{>��$��r`'�������@��F��8����[;�^/�Hb )��i=�<���z�0)�7֚����T�d�Gm�u!�].�^V��#6z�ZdW8�\�h�������:%q���+��"��%��!�82�ou{wx�$�H���N�Ѕ��b]��\`��8�2M,+)*��O[�)��Z'R�h��6c��i��d�ۺ�X�r�άA+�T�����'��]`'G�k�&�8�,�Y���ӒcnL�|��,�hHx�M�1#��svV@�e�����+������U����ߓ0s���W�"��q]x��/F7�&2������TM(����ʳ�5��>̾wOyl1 �B�Ev#�뷛6�*'HX�{�v,_H�	�A�kX��i��&`�>�F���Y���Os��1��ʋ��G7�JB��n�w��I�V��E�Jq��馢"�ō3�w!ͧ���'�F�Tz���%�T*�Q�����Ш?�y�����l�׻�v�6�������Z��|NTD��d�0�^����r��Դ?��U�9���_��\���LΎHO6^���t���`�`�-[W����/���_C ��(s�o���;4�҅�k��(���`k�4&��vU]!W��ԥ�L
��~�}W�U¯\J��D	�M�P��無����'����d��%��Gb�d/O-\�W�|J�Q\�#xP��	�^S%�V�-'/��U��='���0�W	��	ڿ�J��FS!�A�$�`A�ܥrg�/�Q���>'1��6&Bb#΅۔ Ћ؏��8AS>СE����N�u��]���	T8씚:e��&	A�ũ�Q�U��NK$A:�P8J�uq�+$�y��0>�J-�@f]���$mш�k߷�-�bgQ �vꅌ��8��Lk�`3�0���X.�ɀ�9�k�1�;�UC���>��dg���=>�U\'�S��-AF��꺷:k���6�i��L����?+��+Y����Zr�dT�%�y�ۂV�	��}�W����c���{ߘ��;�t�"�ԁ��2)˅C��Ҁ6*�I9�� �p��ԫ��:m-%�0�V�Yh��� Z���kmV��]����G��+�Ȝ�aEv�W6G*6Jȼ���9���u^u��n��5�߯@"�&�I���̏vtP�O�J�*��l&�a��ڎk��w�!Z	b������ϝ?�Yȫ�ö�%xw�3�חr�ԅʧ���A�f����}��zQ�9�l-�x}�菢�b2�a�����v�Ĝ?;@�b��)&�dq�_���W���l�Z�������m������=V�c��X_);�~�lK��m�+o�/sݥ��'��X\������D��&n\�'B�g�h��@�9u��1����Д��S뚙fD���ܦ��"J~/�O�E/�$JҨFD2�T6�{ ��d�;�<�H:,~��Ç���u6`��:0��'���ا7���l������H�A�u��J�X=kw&�� _�M�01f��n�"Lyv�UdȔ]��ZU/+h���q7K���+�m5��!o����]��9������N߾���r����_u���Z��j��Wn+��s�[�A���ד�V���#��H|��5b��<�R�No�
����^�h���ib�&3�����<Fяz�h}d���h��vj�kHCyڕ�����b�}���A�bI���{�:�Uc�'�/rU�Ĳ�o��QBK!�i�n�p�D�y�7L�5m����݌ھ&.\�<K�)������s�쒬h�$�ᣝ4	x}5����c����^�.}��w�8���/rs���96�c}��p�;��o+v����4$�@fL�@�K3�� D%K<y�lg�	k�L~���#�V C��E�L 0���*�s���6A}�` ����$UL�{#�W[]���-��gc'~������l�E�Q��
"�U�G|N�E}�%�\�]��.�O$����U]�������YEӐm�h?��k9�h�WRq	d�E0rLCՙ�p����o޹m�)צ�E�c@ʰ�o]�K�A%�X�c��d)�a��q��@K3�f ����z.Y���_w|/Rؘ��� \QΜ�~(H��L����`7�{�z4f&��9�̕�u�Z|�4�,#{|�O��~+xk���	��׃����Zk�v���aR�ѕa�����۩5r7�oյ�� ����F���#=�)�� Ӹ�%���ОΈfT���Fٲ��*>Ϟ���լ׃�+M��z���SY���9������~�Hm9��p:xy�efp�Tc �N�K���ۋ���&�S?y\��ϋ�M� ���
��q�6j������?c�F��?��[�����L������Ni�I^��g��%��;P�T�?�hv�u�s��!���/�2v�����Cx�E8y��Ɩ:b(��/䒺�mi�2�x��"�Q���@C��X�>�������<._CX�A�*�Ez�{�i��3茇�>�'��vK�&��Dg�k��)��~G�C���x�حj���OgIB:�7�$2q��X�N�l�(Jaټ_ޗ�WM-2ߢ2�;��5���by���Ϟ�'^��Ȳ�e�m����1����d'��ԃD
�����2�d]�rs��q�����<��xW^���͑~
bA1[W���Hg�:�9�4|�͆�M��_�E^�W�Vz�����!/�Оk�Ahr`X�o��N�$m�*��_f	�ǶB�m�0K���YV-�4������L.�9A6�X���08�O���6/�����:���K�>"��Wj'�'�W��fXq�k���~Ҡ�>�ڠ*MW<�}j.W	S���i���!~��:�C��g��e�k��;�ֹ���w��P��L{(y�T�bu�%���"$
a�K���r�$���%�w�j0�� S����/��kq��o<�c��/��
�����tξl����SeS��a��'/��Y�.˭N�����o^HcN��0%��@#Q��>t���
+U��לTv+�@(�U�L�k����REp"��)W<��K7џ(jm��Ǥ�UI�!�^����f�F��kQ0}PC*^�?���U[H��̧�
�����t�=�n"����^�e.�[�����c�.|hOc�$����O_�e�%j�w�M��:I�?�k*EB�l~٣�I�Q^�@et�lʆ��*�]���3�`�+d��pO�BP��;Ts���v[F�����[��� yp�}1�~[��?�{�t���}��zhǏf<A1�1��YrGi���ShrOt�:J�
����_�}�֕�w��w�]+��jA򋡵�:D����g�s��X-5��__N�R��A���	{W�HdN@Y<���3e +����r��1��W����H��;���
�C:.:Z�@�x�{$ �J�#���{>�f��ʇ�O�aG �)�0nEh
6�-�p̴4տ3b�1��ʫ4>�W��$AbL��Jq(ف#X�Jг�Wo���T����FI7M�~ѝ����?\G�?9�G�w�����̍�9�?��'?���;�;ʌ���D�k�ǹ��N�V���5Q��|bv3(j��p��<�Q�Q���#�6�V�֠S	έ���{:�A������ځ�a�}�l��NiyLj��љ:�^+`�M[+GL�O�teK��m��f���0�WY��1��}ʥ,��ݔ#��$z_:Ϙ�u}[��@�E��/���xE��_��f��J�w��Q����l]=��J����m�T0�<"^e��,�#�TE�g1�7����x���+>�y�i&O���Hjtn����Hb���co ������'�����tp�����<7b�g
ʙ6�Wu�0(��c�1s�'7p�dA�HZ�j�	�삻��?xo�'�;-��Ax�e2V,GB��5��㥓o�}�tl��ee���|���C�\1i�4%5i�����[V�M�/*�:�� ��:=7���fE�[;4XT!g��5��,]R��CX{���3fȻ7�P'�J<����e=�9	��xW3�HL��\��Ax��>�9�1�5�P2BmJ6b���n�*��1C�,�qVʹr;�~��\��F�/[{��/C��K`��l����,��r�J�{r�S
uD�>2;Ȕ����L�AXM��sG�0���|p+��AP-¦>�~�Y��Fپ�x6J	��#H
���
H�b:��k��0�閹tE;�rxٕ� �������2���\�û S�Ӳ�������b�g(~������6ic�LJx�{滛Iox��Td�`�qYI�ÿ���G����)����L^OG�%Z/t���� "0 �گdE{8{�o��~;'6�;�kͮ���D�9�*�jZDSⱚ��˴�'ށ��|4��[��p���r|GB��A�=c~ t_ ��M�X-�.�9?I^݀10��3��ht� Q%��F6�	/B�_���Ы�mOj�<�eta�(D�8�k��Q��D[�������>R�:�Z˾�À���7mV�g�_����jE�N9%�%Q`s#ߊy����8?��xu��X��&\���-k�4^H��0V[�=K6��ȅFS�YУ��h�a �dP���K�A�|�T�o� �)v��E����BX�p��NWi���� �Y��
��2W��զ7�i�����u�3��%�#�rjO�N$��/�^q<ֈu���x�P&�@#��&_��"8��D���-�@����e�u^��E6C�k˲UR�i�fq�y��˦_����w ��4(�s_��]G#bw;+�d��T_!h�t�a��`n=�3����sܿ_8\�cT'������'�EA��np���J�&93ٱ~K���'���Y_�Z��Q�IUevI"����a��6R| ���%]9�����ȉ��@�]-C���E��j�r���uyL�)*%<T(|��i�A����n_^�­�*���]u�蛫��G��]	����j���eM���KW���M��Q	��\���A�`�kd,�{pC��~���9�!(���=\!NAZa�Y��8#�ҳ\�d�P�խI�����Po���va��V����1� �}'�*[�,�*V�)���bz�a�Id���b*��dLe_���;� ��|�z��������3�*4�	oy�~��z�+|2t���<��C`�{��wv�PDƔ>By��	rqB�OD��qz��*���7�`.�o��fp�m�I�Os��s��h`�gT������бz�\�!f	$��*��Z],����L��T��Ab�{8�(��$ 䭕����.�'������1���1?�S�ӾE-�����v�wxm�y�C=�5��qa���;� o����ĔQ�a=�ř��K�]O�ʖ8�,�6_�aX��oޗ�2ƹ��eR�xB��J�z	��ڜy�?R�"�3�om,XFh�_$d��bi�L�{I|�ur/<��T�)��_M�E
�{�i���lBSk�D�p�0�b�y�����6��a�i!�b��A�1�[<�n�L���>j���@�z�y�0�>��F�{d\d��J�^:!���-<i�
�p��ͅ���3W+�{�j�jL@�Z*��4��E������r���5�ͤ�.W�2���B>�J'�xd������'�N��j�ٍm�۲�	W��%vF����I�=����}۩������a~$�4��"�]e��s
�����Ju�\�:�pء�P��.���
�腳 N�i4
��ޚ%��i��.������ĩ�X���)��}i�xU�)�d�`�*M�Y�{S	�1QV��z���Yiɉ�-��Nzx(^���%�� ��`q�Z�~�a�D��T��Z�G�a(���?(�����˘Jݵ���c	T^��7�9!R���>�	{$�2S,�Z��a�Ԛߤ�m.���<��:J�bL�1XJ��7��ជ+}Q�^h�B���枾�3*�R�Z��{G�NNE�z*w�����ɼzjV���|�e4͹�%c,-ƃ;��c�ܠ���7K���LY	�Gx���s�0�7���j���z�L��@T^��֮����5]�鐋2H�T�9�+��t������������s�OX�]I���w���������~��ɗn��W��	]
E;m;m�oREZɑ�Ң��y��u�I��LMv�jxelG;' ���Ϸ{�Ğ*�jXQu`" ���g8�a姿������\�X(�:��_;�Y�#�֎����"/7�/s
B�c4���Wm��4j�(�6�Hr�ٶ;�Z]!Qʫ!�gɒ~Q�{{C`�`���"�Ds��QmDf������޺EA�/�F�7~f���e��ґ������wS����_��(~9��D� ���ذ[�ed�ś��,TL���A����l�3n�H�'i����dv�(7��	@˱�Ӱ��{YW'�V��P�&	�Oo�������"�.||O1���ڂx��4a��v�������BYCYi�/�΅���M:�%Ơ��S(~��
'��~Hjj��RXhtH�E�7�r�J�S��b��~��W����o��{Pf�Wsb̿�糣��L�[��*G��8Ҳ�1�փ��"�Zq�	�:�8�/� ܷ|�AO@[҇�	m�_J��Hɧ4�O��V��2_~䖸�ˈl�D:x��p�|*��{�=7vއ���
���×�z��l���'��kbt�HG�K�퐏|&h���1���h����xg܉��6�$?c��ST"w����غ�����À��o�x�=�?Epf����O8�z}�E��nt-VǪ؅n(�jsN��qm����q^��xO��?��AWH>֙�����ɷ>@Sa�`T��b\nB��H��	B;��඄�q���)�����C������v-<N�QE�ކ�/Q9P��b�����IP��э��6��q9�c�N��}����v��9��c,��0��Q��|Y��&��]���I��q�S���;Gt�����)��)�F��ZwX(��~�lqe�M������4=7_|M�lԜ^�ek@��g���?,	��1g��7���S?���5j�?�����0�[�;Y�sNn��$���5�h��%��m!��e`�t���/�n�0y��EZV��S��y
�7W�\��>IY�ݐQ��x�fv�-���Ip��F ���)O��S2�ʣnώ��D�D���C�N�q�͇5^�I�4�fL��/�C�UV���H��W�4B8}����R2�~CT�����Gx�.^�F�s���웺ϝ�j����/}����~Vj���P7"yݟ{\�u���e܆!��'�ɚ��!}/�	�k�"a���J)�Ɖ�!�\���<��P��wo!	��	�h3�RT�xN��{9����}���NN���/����\�'65c+�LD��Q6`6<XA��,��_��.T��la�Q��P&�R�b�������uC�gʻ��S$����O���I�̋�o�#k����`�V5�r�!�b��մ�Ae�'�~YB��ک��Ӿ]��?�(�E:��-��uÌ�bL�����=�@ؤ�\V濔�|c.ǭms��n�F��swZ�C��P_4�+@玎\��U�K��'��"�uA#�����L7�����]��M^��{x#�P���0<������s1���Ox��1�x��r�]'���7�J`�װ�lp�wܦ�������][�3����t>W�}ف��͗��@��2�UR\����W_��\P��Z9%�!����ӄ[�%rAP��3R<]�#5�L�Gy�)�38��$jG�����	�5�m�a��7����
�9��p��`�,tym�<tڭ�l!߿���B.�K�[_<��K��r�R�h��ށ����:�>"Ϙ�\X�zy��ߡ\���a���Pu�T���>�-�8♄C��;]�RW|p�a�)�v�}ũ����l���Ia�$|�`��L򮘞�##�7g��nxD���x��9n�J�Nit�t�����<�S����*�>���}��[��	�
��jݼ��Yz?��K�	MX�'f�[+Ko��5Z�<�Ἇ/��Od��ݖ��9�3��Ubd�]KB2nn�F��<i^��Ƕ��a,aU�x�46ٱZ ̇�;�L�e64��H����/�4-T�ߺC_܁`��e�����Q~�?y��X-�YNCg�$�)s�\q���uw`�@fӛ?�҉q.�B0F,Xe�}+.�Wc�}g�!��ԅG� �e8{,?���|�c����(��eJyb"oj�wl�,�ꣃ+���2O�����<n��� wY|@AQ��&��n���?���J��g�yIߤ@�*�Fn_v1!���y��|��1���5+B�E����g��UUA'��}�4���m.�x�\��3m�U*��~�T>_'�v��] �5�l�!�p!�2�7@�W��͜(ބ��U��`���?�sN-Pk¢<�M������Ԭu���%r� Au[��=[̀��1���wv��e��hK��6	��~��!n�;ej��IfS9��Y(���]E�D�o<
���TY��ҽ��tx[
Ç��O���N��O^,KJ�������ӻΙP��bq�C(��T�4Sec��=���p~�|�Y�=>��A�I+F��x骷�%0���g���҉{�?�G�F�b�j�8u�X 8H�Z��(�
�֡�z��C/����Ex�bf�����t��Pyo!�ʶ� 6��D�2�*u�7��& 
���֤nrƤ~�L�Ͷ���S���s����_���Tю��r��&G�
��f��o�H��`�~2�:��LI/�m$�XP�ڇ��:��R�C�ޏ�)�P�X0țF�{(��\ל�N�i��pxv�m�,|��j�F���%���=���Dp�v?p[�9R]C9����H�LYZ�lC�����"/��,�#�k7M�V�ї�����
� ��\��`���W���Y^(V�e%Հ���n�� 0�S�� ��-�;�ȹ���(M�����jG�6�G�{�т�)���)@?q��f
�<��R 
/�Yp9�y\��a~���竌�<ه�lQ��i�FOB����w�/g2�R�O��������*&����AQ�Ȯ��FϷ]dR�����N��퇩{3g�.,�F���н��k�l{����ߨ���3Ʋ|��`&w�e��]u�v��}�.�,�V8�QC��R<�o��*��i�D3Y��%UD�i0��2K�O��(*'��f�@������J&;�9��lF޲(����ZN�~������}����a��>�� j�}���h�-^���H�5��lB�^�Q�t�WU�1,�O�b���v����/����8���J���n-."������ �P��j�7B��܍����Te�qb�=��ɥ�&��mvl_V�Eq����ǽ9}���H���7_��.�GVQU\��&���%m��1M�;ev�.خJ���@W�n�)X[�荃:II��V}r���nE!���^×��iKY�Fm5eBļ��8l���� �c�%���]ԡ�u)�e�b[|^�X|�Ɨ���G�j��E�4���6��sߏm*����	f�)�1��
@�a�[�ߙ!��0u�G��� l.�f�ȟ��tyRGuVF��x�tEB�x�� � 4ҍJIK�kz�[�,��1��&_��# �@D���w�V�Di�"�r���6��>Z��J����'Y���#De�G�P�[����Q�U���ru�#�j�c��Y���fW�,�p�.�O��1n�3�O��xWn\W�zA}���F�~��Y�I���U�F=���]�ĵA8w�o�ǈ�+��Ž��k��ZT�7ж�Їյ���+�>̖Z�t]� �8V�����õ�ژv!�$����^x�jH �nȦ d4�������[���8�4&���F����=l(UK'���Klu��E���Y��B�W	Mk
3'^��V��^�:�~V�zʒ��$v삏A��&zF�Y%�:�q�N��
�F�N�,������'<�!�=��N)g���=��7��vf�?�Y��|�F�D�e�@������Aq�g�\< ڣ�|'�k�����N �^�g6?�3�u�*�9���(����%�L�蕤/��a�c3,�����^�)��������d�������u�%Xq:�9OV�awMp,M��^g%�.eT�yg�ñ�!��k���YX�x�,�>����{��[�2�[�d����F?�T�6���Q��z��#т��LG�$�7t���T�=�SF�3�U:F`vg�9B#WĈ��v<�j�$�܆��{z� ?Ē��c���#�p�S˱X��7�ހ�Y���xE������}����ʡ��on��	�̾����L�o�kvci�%��t�����m`ɞ�0V�tXmȥ��tH��t&�w:�&���B�2�5�ш>4��,�mޕ�2s�?������Yj萌�{Y0�4х�