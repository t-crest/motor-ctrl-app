��/  i�ί�JO��«�ȹ� Tbp�o��2H�F�ڨ����6�ԢfI�>to$A*�m�#s>m��cyL���R���kYD�+fl��bH����t2����3H�^�qlvDӡ�v�Į�5���FS-�ތ'�s����>V 1D^-���3��µ݂E�^��<�J	9�yI۴�:Sހ?�!��mbH3.��^;�b1�A��Y�Ǹڢ�n��0-��$I-|aqa��w��B����mk���W"�l1�c�������!R.��)'�������R�Uݨ<힡P�����WS�vR���OS���e?q'����gKS���-o��Nr�K�,E���-��ufm�#�2�i�$ai�%��2贩�� O�~��|�C!d|̲K�Z�8J�MQ!t(!A��"�,���C|Ùp��ŉZ�Lgz[���z�(��V�-����Gt���Z/��tb�{sl<-z��±�WE^0?����ol_�mW��ߔ�G6�ht�,Xф�su�	��i������ʃ�Mb�])�_���Y@e䟮WK�Ym�M`�%<�杫��Q��0+j�7�Z��򃖎ݒ}�A��w �������r�Ѩ�(hQ$��Ņ|������y�p#�.���1`rɟ��K�!Հa/l�i�����Q��2��|)|9�,{�н���巂��ob��t�8�݌rM�XT-��Z�-�JPpP��\��]��"��;.�=�0	��+��䒐�7�jV	U��6�x�oAWAy	�[���P{SLV���s�B��4�����.ۂ*^+�+ �x}��ě����-G��w��m�%I/�"Lc<K☰~�QL�Żﻍ*����t�.󺿎̺0B�H_u��OuUn"���x��Nt����ڙ�3����U�n�f��U؝�XB��e�`��W1�6d�� �b9�],�'��1%�Lq�������J��Y�/#��_����#�s(r6|�ع��v�����
��|x-������kң�ݛA�GO��\'�00�~��8��t�S\i�x���*�Sl�1$��Lzɝ�Ԍ�x�����:4������8 �r�3��T�ҍ��A�Ń�����؃"å"��7B/򲙒��c�7�ܛ4.���^�����Q��d�`�Ա�T	M�eM�0χ�h�f����M��~pЫ�+]}�F���5�h1S$���m|͋\ч"�g����5�1�NO�u�lȆ8�����U&���x��n9!%�[��j���`[�1�3���!R��l�1��9n�8�}��{�DqhF&n�xa�ao����3��o�>Κ��C��^�.���KL6���U=��V�Ăd���H~��<�|��dy�h[|���@:�{�(���G����� ȶm̛΂�?fQ�����G;:���_4��tc����JI(r/z0���?D��i�}������1���y��.�L�;�)��.d!��jj�)&{�u<�[7�}v��Ͱk�E�L��*��,z�M_�Ft�\��W[��y1
����I�����9J�)���}�ȭ�R�/ǟ<������u֑p���&��y�D�x���kg=�rh''� �X�����P�Ġ���;��_�:��K:�T5�l9��@C���8��p��K�`�	�'^��Y���@<���I����$��9e1�і�K������W���������S��t1�v�j�q����cHt��'B����-H��Z��#�90�9L|�}qT_h�=LEAr=	��&vA`��>0K��T!Op�������u�l��1_buQ��j�s��uI�ؙ�cnYf�,}������ 7#�9'AB`��BW�����������R�����חػ$�ڛP;����_�y-��W�k�Ӊ�DW�t�\J�A�ÿs=��$ Ǭ�*&��r�R�Fо�u/�Q�Q�6$S�3�G����w���������xp"ɬ�����uc���3���p�]:*���89����֬�AT��6B�y^P;���e�ts���a��v܀׫���d�rRM�
�"b�v��p^�����&%Y�w=o��ڙQ��0��Q�xe�����G��\OuT@�1daA#���W(r�o��#R����[<ʎXɦX�u��!�q
��DDf��2R�l?m���ni#	��y\�v��츬 Lc=��X��
�
Q^�6��Ԍ暆�(�5�U��$ꑮ��]���.oWL��!�t79*�+���6EB�����2xxa,�4���VƊӂ�78��M2�rѿ���+���Mno��3r��X�2�ȤXl�����#)YH�|��k[��%���,�����uR�M�����"E��ݍ�{9�A�j�eS���[h�PN����Z��2�8�	�2G���=�A<3K�g��g >�L�s{Txe��i:��T�4�xK���'D����x��+b�>b���G�ջ�p}�����ї;����O؋��~��x��?�2�*�9y���~P������,��ߍ�~e�u�=������V���D;$�����]�jO��oα��i�<_��M�b\r�h��_�����2�UgHfmv����FUڐ�	��ϊ�'S%��A�.1�1�C�PuAZ�ۺۨt��?�͇�� ?`�֎����O|�.��b��	�/UI�e;4���VPE:j[��,&Uhe���ؖ�|5�Oq��[�ǰ��@:��B475�dA�J�8���v���Q�����X�PSm0ԙt�<���o0��L � ^������"+wf�|v�����'<oRYB�&M=2� �dȄ��-@�:� ,�R!���,�R^�ר[���=?��!-���,�Ԓ��H����i��)^�3e�7�n�0/F�;�Gd!�� c�{7��w�m���Ŕ�=HK-#ڹ8_��"�p���~?"�bj@g)�;�l����wSp�/闐��y�D �(�/�Nz�I�Q^ua��2��H�+0=(��a�{��5��.�Ȣ�K���{X r�nѤ{3'=<0<y��׈�J�>���/��D�5n�몡��/Ӡ�R)�U�%�p�;wQ�_']N���xV��I\�tSV[Ύ	܄����]�� ����Pw{��u�LнvJL�ǭ r�t ��
��3)�\#��2Lf�EÐ�9��tS&6���I/�aF`d/�NL��C�=�kl*yQ8:��?���Y�/�&.u\���)r���@�E	`[��*�w��+2je������h+�u�a��~���7�J�e>N]X׽W��>l�����D��A5v��y�)�7��*��3�j�qx$�rZ��*�k�R����s�8�0����������|�ЊD�n�1�^��x�G���ɳ��(>�#���p1n�	ǖ�����lu���ū& 5�?�x�j�T��wxy�9�Y݅.�o\���q56��G����B�U�����0�4�����ɭ	�'���nAE���i���;<������<$�	 c*��L�kQ ��<~�������_�屋��N�n`]�N�g��1�P��G5VN*�F�VsVqok���ra d�WDnsgK4��T#^���l��0�e��goՓ����ˎGHܖ1PD|��ˊ��F��h�k�N�m��I�����]s~D�1�ݻ�y���˃o��zl,�3���Ȋ��ǑB9�.�	�+Z��g|&�� ��pk�/A9�w��sD��<�g�1̇}�,e�?Op�Q��y�=Ӟ�:�C�n�l��k��.�+вWns¢P^(Z�PF:x�S���dڂ3t6���.Jxt6���:�h#A�|���`_�K�����/�+��8����t/rrHǊ��h9Yn�m+$Hb�өQf�:*W4�?(�S�K�Hǿ#E��=�BFpq�� ;d=.؊��Y{��2'O �Ǒ_�B��/6u,�$�B��������r+WM�l(P?6b�D�܄��[�@��K;*2L��3�f8���R�l�(N �x�!�#bӠP��v���
2J�<����:�}����p,K���	u�a�+��J�� 2C\I�	?%��b��qMN&�ԽM�H`[
�c���}8{�� ! �˗.
���F�Tʐ�b(���h�m�|�/�8jK&�t��_�sײ�u�H��Z����x/��(Y.p�~����V��� �:w�`Ȳ���%���6�&�F�6�Uav�Ӈr�Z����Uo��#�b�ȶ�yDn�D��N�3A�[�^�_[!g�DՔ��&mP���RYL2�����D��h����ޒ�Z*�aU>��Y���r`t�th��U�@�v�=ZjC�Im�Mu~E�KR4�n��
9��{4��)`~��p?�k|��Y� Ѥ	�+*�?a���E��Xr%e�����z: ���ilDa��/,��u�0eX�F�!�X�����2h���([����Ѽ��(���D�ACӥ�n)wfd��7 �w�4�L$+�%�����RKb�'L�F:�p6x��V$0Ui���c�U$��r}�@<��p��Q��_oN �ꛨ��m?�'��gv�U�fK[�� Nv�`e<,��@��JN��?Ӷg;�*�@ئ.�g�xqK��Io����(U�u�Dd5���c�~1�nw����ma
)���^k��S�Z����C(��Ћ^���@�Z��$Dm���&�����_F��[�e��j��<�:q���\���p��"��.�b�(^���k�=0��en�C���ȔӲ� ��`�O���o'g,�"�|��S畑��փ,]Q�u�|�����]��i�r���4�9	�����Cˎ�y���^O�u���yX?~���Rr���#IR�n�w:4��ͧ�����	��1C�8lGٛ�U\2B���'HNY�FVo
�I�����v�ҺtcA>_WO"O�ER�ޚI��<��$K����U0��]���D&�J�]�����Fkn�J��Z�9����這�{Q4c�����vK��#T����җr발9��@uK(,��Rb��ه�lnP	u�S�?'��km��IS1�,΍�[�u"u぀��Lu�$����~�.��e�yp��a���������l���uS������kMBD5�۔�/�'���!`�"a5.c����vl4��ȁv�IK+)>���C&���^σ� ����n��B��٦��lW�}�PtřN,|>�CQ�'J_�����A�[����{�c>7"Qi��տ�9�%�h���9;8A�D>�ߘ��z�M���*(�E��J��W�q˼� �f;�Vuy�_�c�'V��	��Rr* @lw��%g�Y���J�2/Z���*G��DEq���c����LV�?3`���|�揁YD��Ϙ�`x�1 t�m��ބU)j��s]P���sk�H�������B7&�sǼ�Atfq���UH��E�k˹�W�#��GKg)P�3��R�>��G�������(О��/�\�W9�w��_cT a���t>a]��_��]y�.����8�!|�A�k�����v�^N]�-��޲՞ѺK<���%�2&�`�*����W���v#��}�~�sFd�0$!>�cȏ32#�	�,w��	އ��!|J6���ŀ��^�\��+"n��V��đL�e�%�N�`.�㶚BW��c��z0�=�u�mb[Ȃ�O�%$kض�������&�ݥ|��_�'�`r��e �"��/�CU��M�7��AQ��Jt��+��kn�t���_M�nf�6��X�4/>����t��PD�ި�o~�q��c��ɜ2'��.���I`�>�v.�E�8Y9���"5��J5�g��F�3}��g�?�V�pP!�tYT�t[<.i��z
�	
�	� ��o�kN�ɚ!7��gpR����~��j�Dhj����u�(���^أ�L�� 1"�]�n���UV���M}��J6�iE�M/�?٧v��AUc�W��%e2���/'e12t,GH��X�JG9�I��)g^�n��D6իn������54U'����q>Y�CM����a�<֤�_��Ԓ�,�߈���W,C�T�JYY��^�?;�c��	�Kֵ��N��(?�K7���>(Cbѥg.���v�.E��E �|���٫s �=
˗W4F��'I����+D�"��aWs�h���to�T�|=s�=: ��qd���7�,���K�? �.{��l>xI�p7L$z�~�#q;��}!���%֕���Ak���'vE6x_�U�rc}��z���S[��ϼ['��R�drr��B�aZ��Uģ�ޘ�s�}-��@��`<���w?.�'>�2'��b�:cE��W�_B�`���S'��6˭�o>��1p�ů�g�Q⪯V�E�euɰ�[�t�՜�1T�A`;��,�h������[�҅Ɨ�G_��4 ���L���/��5��>���{�bÝ:�X)m����e�
��7�'�(����7��(`�)-�,Tśݕ���ᚅ��K˕�f�)I-T�p�d�m��� �gJ��6�(�\��>�+'��z)P-nb��{���|dL:Q�^8�I������>e�c�j{��0Z�-P��+�H���(���x(� �+��$�����PV�"�9A�z�ʂ��;�!S�,F�c*X[�T�C�K��W����6
9�nJ���o����	���E�%���3V�!X:��5u��v_��Ĕ�f������>�\�iȊ/#r�}����w����黁���Y�k�_�t�ϴ�V�
re?h
q�Gf��ېb�����"���wu��bq��ǈWy�X6|<�8��'T�rK���FE�nc�+p��y)<�L6���)����6���1��a�$�<�/Ph�!	�9��hW+?)�h��5�������W���A�����X1ҁ�AL���L$B_���o��`ec�^b��ZY�m_&Y8� ����s�!}��g�ihZ|�7W��@k�`�ҳDA	����0d����OhV���@� ��ѱ���rXG.C	�&͑B��#^���WP��}#�y��N0viҸ8x}>��&P^mg���6��f��d�g!�u����{�*]Ɍ��0Q��L�����\d1�2���[UL�"t�|�t��DL�T���Pj�RI�;C1�0�q&���뙫r΅A�����X�ۘ	Y!4��y���Z�8Ў@�tFE�rY��;��� jy~�pL^�q���1i|��8�Vb6Km]c^�}�MY��I ;�"����<O�m�t:�����gP�����0E��C�s"��C�OfĴV�9(�G)o�b�"��;����#9�(_���=(�����s#���o���i��'�u��Ȭ��h��࿖�*���e���Dwa:�{�~�P��ff�"u�"L`��� ~`��3�����3I)��������hn��|pu�̱&`(C/���rG���"&_�&N�z �dvi�`�0<A�kMդ|>7i�C
�9���ys�A��}Z`=��g���U�"V�P������Cz�ăAM�-.����˯��~�t��0��LR��V�\Jd�|F:��Tb|�FS�l����E�& 9	��*��c��{b�U]gt��w$h���Q��1�8䝸�mV;�1�JR��>*��޵��J?%~6����]���m!%�C>��u�����W�� _xA��h�(#RH��c!%��!� IL�8_�������hT 2.c�u$�s5v��S�q���g/{-l%�̶����FB5��1�]5��n�J@ �fǴ�\��1�s�JX����P[���s۬��k�R�Q�H���p}�f�R���7&J��Q+��L����T�������� 56R����D�Y�y<Iawpy~M�:S�[5у޻&�N�<��*<U������D6nh m?�Q���7Io�5�dN�c�IֽP�����w��poB��Ԝ���Y)�>�a��Y~;9����a��Q���&C4���9�B���D䃅��,����ȸ;=>�lx�[(�ojE>'rԩf��zz@�5�����-��v��,�,���˰�"Z�W�a��]�j,Zʃs���P]�����:���W��`WD�]��S�E*I5.�xҽ�m�*������C-�fV���F�7`�k�b7+7:�kk����?Ȼ�MZ�z��|`����d?�,cR��(S�݊ڔ�Ҥة�w�L{��O�?n-*r����.��e��d4�v��mCA/�h��E�P�8C��.�p��e9"�L�֍�y�}V�~�BS.7���j�)�VH~]I�g��^Rh���H}�<9@g�լ���q�m���H���-/��^�X����7_:�o���wO�F͎J��.?Y�	(��'�o�Qm��D(�9Co�I6h���
�U!� H�x���[l��L�{�Ic�1Cb�lƍ����	h�6�⦹.��tNWP�