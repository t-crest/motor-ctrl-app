��/  *�>�K@^�e� � C� �ѩ��]�G�������L)y0}���$�ﱀ�]���0�(j��U	SM�2���c �q����B`aݿ\��bt���y6�Dɷ`�<."[�8�$cl*���3C����W���*���8�c)��ܾߊ]�9%{������K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<��G�y�F�W�0��c�X) /�Z�I�.�[@Za-�I��=Qg\��՘V;$9��6Hon���8�;�c��s��Kԣ�O �e#���:���'��qK�EH�9T�9�W80n��*G!e�[���������B��s>��h�K���?UR&�MDG���g>�����{{���P���Qc̬,���	I�e�01�9�ô���,�~~.�_��h��@o��g�9�b�k/gl��Ou �r�"l�4�x�NQ�����o�u��
+,0O�>��Ͼ1W+NdAA�r@�R�@�%���&b��%v�{̗�);b��~:���6���&�R��>��&>ؼ����O�p����{��yp��Tv5���}��vãҰԬtX��,0�N�86>�Nݭa@�Ȑ�v�ܥT/�d0�*E�q[�~�7��Ws��Q�W�,>���*!�n�k�'��&�4ǎ0�!��G�?�S])D��|$�e�
p(���|��46��f�>�ʨ�͊�����70MGd�!�aw�=�?3��p�:��R"������U��H>>��ڙ�b�l�wi<-�7�&qF�-����sO�Xl)�TW5"����A��ၡ���Y��:�A�^nAQ�������#@Ɛ��u�:Yӫ�?{ҁfY��S5XO~�_H�,=��\½AM�C���u�Yw��A2���~A��w�`�kZ0���8�۝,�|��v�����s��JW��8蓃$���?��>}���<�9��z�����?
��\�G�3����x��X��A�2P�$�w9��$z$�k�����W:c��<|��F-�q)�y���pI��_+o�Ў�@��|��4`��Q�����9��4�Υ����<�L)Y��������"�����OP�dx���]a������~�N�v�����X���_�� r|8�����r��<xA}���^�a�
U�\
4��+����1�b���E%�e�C_Hh5@�'e N(4��'�k�l�㺜���a���\�ϢjReטPw!��KJ����]�	��S�H�FGl.�I�e��z���4J�qmBc�S��A��D�g��1ZidE�$���ի�0���LQӺ�)�h�m���p��+Ru��OJ�vjCԊ\GR`u�p��E=���Wˍ�`�CҤ%Q�M��-�^W��i��<&/���&D�I��0*�X�'[�Ӣ���pm�=�1�#GeSN�P��E|}���O-u8:�0['��
�S�t�P{�?
7�n�M�h�E���ḷ7��y�6YuU:]�z�R���}.. �b��$��\�rFR>_�ō\��ԙ�zO�gr	��4��.:�Bh/0<��D�D�E�4��XKc���.E��/�2j�}�}/ɩ06��}��	��td2��2ׂ�$Ĕ�g��}+u`q�)]��3Uj(��_غtS�`��m��:�@V_�`bAK]�\>I�yO��׌Bpi�dd�K{3�3(����h˔d.W=�_*�lY����׭�|�z����h"�4c�X1C�+��r�=pD�E���ă�)��Qu�3A���_e�Q>��>����W(-�v�v�K�c�tc�:����9`�2�j�cu�ղ��>����2T�.Y��X�Ѝ]����Q.&XN�{c��<`�?��V@���H{o��'�3��F��@Q������|�S��%�H	c�6{Z<�`�_�MB�8s
�bG%�j��/�$�Q��̢q�����_�#��o�r�l(��LN�K>�: �q\��h+jw1�Y\�k~Y�#�����>њ^����tm֤���6L))��X�Rꜝ�L'S�nH���}�_�HN���Plû�n�#�A3c�n7�驖ΎI-�"%OÂ���(e��* J72��R[����e� Igc���
͉�q�ׂBʣ�ʿ�!Н4�W]��t&�9�O���-rRa�[��|@T��F���`Tc�6_ː7l�����̼�⊪�[��7Xܜ��2$2Ni��1SҶ@V���@?����b�?�`V6�<�}_�cv�G������ }#�o%��,�+�NMc�6�x^�����7�	9#��f6��)��tَ����OG0���� ��\/.ߚ���зl�-MDg��$'�k ��HU��5Jg)@�e�2�z�Rt��h�Q5l��"��=*�����! J���iߞ#�.�X�$�V��<h�`�����WE�j�>7^v_��)x�u���gV�?���2	�!�"k�~���h�;X��U��a��(�ە�D�u��:ɏ�ߑ�%�עX�ɔ�P����}ۃ�4��(J/٦��0(#��
E��;-:�L]�U?��$���]ѓ�s���"N�/�B�aRj��6�8־��y���ƙI׸-B��/=�`³th֙o«��������*`�����8�J� ����X3��Ļ�����1`	��K_�҉&��u"H5�B�ND��b,���ЛR��[`~�͡���=	E�-D���R5h�?���?҃����O#�ur�U(���*tk�o������81�&Wcq�o��cT��YA�6�>���iuw��@���踽Z�S�A��Qs\�,eO�:N�|e]�: ���$T�����@P�f��q�oD����`��[B3��H���$E����$�]�G��'d�6>Ƈy���z��O�x����Q/�©A�*�������Ƃe��)M��/Y� ��Y��K���k�,��}�Ɉ���cG��O������_!	s33=��u���+{�*��PS�>l�ys����*_^Ц�� ��r�4���4�/���7V�2�|�����o
��}����Ljc��Q�m�x�*��:2��FZ��j�B ;�]H��똊:��A�p��ő}��-X��?L�ɶPw�ȕ���#oAJ=�Vf?ՠ�Ja'l+�\Ջ�l�կ`/]2IMZL���#h�T�p�f�^���1�_���Po{_�f��� C$wD�>��k����N��O
�j
��\C���"��5 ��=rU���X�zx���(���?߯ɣ)��LU�3Va!Dk��'F2�r>�����؜(-���(�R��ۙ�	���7�G
1v��Si�q�����!�O��4��z���aNˆ濅Q�X��zîN1����//��7OJ��d�� @��3F$t���R����+�$"n���>[�� 5R�����_��(;øM�)�0�$T&1��d����wN�Ƭ���US~r"����[[����M�R慷�T]u;���w�e�DG\�:Iߺ�_�ʌ�����4�V�m�������c!��6�hUq�P�?�����xd�A��Vb�i��m�n ������k�g k����[Ϟ෴+%