��/  �r���TB�EL�+���iŒu+o�4Y��0��Q@f�q8�="q��[������x��x�Eb�V��g����eں���G�퓝�{��<6x���TH2 '�C�x������'�D�� 2-����d��v�ӱ��E�� :��V)H[D�l�� ��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!����ıL	���dG׉:�v�&7^ș��+�W1���_� ��Paj�u5�����Q��ߝN!(��a�:I�(�w`!A���t,�L��Jpm�I-N=99N'���+L��T��	���u��i�؜Օ"���i����U�|�6`���')<��x�-�xF��ș���<*	�m$)O���K4��	tצ�H� Ӑ�&���e�n�z�a[%�,*�g�F�*U��=w>�qO�9���p��W��)6���TlyfG��'y��٫ԋ~���e�(�&`B.>T�o�ɮB�**~Vq�5��}K��� 2!�j�o�� ՚�`:m!�|�,�Ν��O�g��"3c�1���H�ُ��Ha}I�V'��/��y�w��Y�J$)`�%A������UέD��ɕ�pWE�3:𢡊��+��3��4�y$�:1��H}_�j�0֚+J��.�;,�}�e-�@��e�\��Z=&h"��r��B�o��F����fVY���-ԉ�Ё	�����,�ݭ�F��f �CN�&2��mU���� ��_�}$�O��������8�g|�g:����rʼ��!U2I	#;��0�=!�l�>t�f�F������uЧM� ��5���!*�Fw0�>���V ��ptL,��m�υ�;��?v��q#N�l���o-�z��!��32�K�WɃ�Wƭ���y�n��*�C��ωw���s݆�h^��B��}�4^eabh�+ʴ�EQ�+���p�@���T�9�`�r�q�>�w.!���$]ug�������.���ʆ����%'z���/w8�W�>o8��ya�ن_2��������neI1|Y����7j�ڹ'F�Ќ�T��YD!:�D��J�&��i��NI�o�uY�ցX%�KUXw�~*P%3�Ϯ�)�r�g�z����M�僮�n��]�F��������q.�FR��9a��8Uv[�A�y�'�=\+}�(�dhKf�e��/�-�<o?v��~�ȗ�m��n�����|CGH���g�sX�O��C��k�;D۵���
&�*�Y���#D	 S�u:�BٔD�ɵr;���a�?Y�ެ9�qP�r%1XԤ������0���/���:�8\9��<;�)�{hQc������p�Z���Z��w�Ԧ�!��Ֆd���[��L���n��E7G-�����/<�-�h��@mWCs�2�A�G�I� ��ʵ�: -#E܄�I[x���>�^�q3��SH@)�q�IY�b��x!T��x����8�U&�?��dG�f�"�t�A�T1�6���*�3k|������6�{��8�]ώx�8W��	�6/Ok�5�A�����*>��w��Xh1�����'�ĺ�mO�QFc����A7mhxߨ����<��\I��/o<��=��)��f��Xdv��)A�� 	�-��U3��I�(N�u{5�{�(͊o�����o��Wj��7J,Do�|�7@~��:�)���j���j8絝.[��,.ۙ��E5��J�=zǊ�M�%�����3X�e�^OIeZi�+�S�B��Ӿk�Ý�.��G��K��A�]��B����#��'��\�B*����:�o�Ǿ����G��a`��4T�3t����7*��0L������9 ���S����u�naTlxI�챋�d��N�򑸼��8_�ųţc��\�y�Fo��
-��_0�W������D$�"V������<E4W<t��O���|��CbzW�N�Őj���]>��U�z��C���
�<Ic�JLP�Ӥ��c)�l�~nf Ǹ�,�J�Z�-	wd%"����6��+��"?��)TT�<Pc���)�[OL��4N�/o�C6��'��(��^r�����Sm$l
�q=2�S��=P�~Roiu��p��%��~p)̳l�t��|=�*���zp���� $J?5ש��G��4��h���~H'm@��4��bVXӽǩ!��}���E{�_i���Ua��o����򽧀cE�3�
(�ǼJ� �z�r;��3S��h��z�Y���.��Ui_�tob�K�ݰAp��/N�Mu1#�57�;8����8�[�w�*O%�D���>�w]ӈ����"<8���f<Df?��o��HƒM����T6���g�҃v�)������|c<�ыF� �7rxCZ�ރ%E�/�H�>�����c�(,���V�dF����ԫbʍ82+���hm?�X?���N^��"�����]��� �S��!�E8,<t6���\�{��<���^�$�<��4!��p�a��;�Y��P���(�l$<J@�r߀K+0]J{��u��nP������o�t��g�s��f�?�@V���-z�q�v%S���ؙ�����ơ^TdT߅�9��_��߯�n~��~�Vjґ�||�۝�(�0�~y�[��4� �)3���G'�	Դ����"�k���b��h�|A��I�G��h����ƇS�4�@��M�t[�q��7���'��)؄��@�Ĉ����T�[��R���Gݴ��?�Tc"B�1$}u�V��.pp��Ԣ��+	m.��}�f��c�6��5G@�S�b�ר˞xЫXB�uBC��,�x-IGQ5�1�� ���s����^�6(E��~_��g\��2�.�k���꼈����t�{��f�ܪ"D��<v���->,l0`ӟ�����ு����kʅ_z���EB��o�tM  <JFP��&�b:��=v�����4�P4e�Uz4:���)�2~�?�4�`��:/N>P��q��)+T�A��I�����j����\�A{�����ܴ��U��P[�Q�*r\^N���w��Fe�@�]:Ҋ4��ǧn�^p�]�Sgm�4�ͷ���]�M