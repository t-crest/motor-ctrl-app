��/  h$�p�̦qQ���u��].:���.���l�v�<~���)�z�6t��6�6�R��@1����3uk�R�`(���������FKv�f^"�	�OdB�6�l3 �vȌ����/L�7����zBR�yʑY;l��n1&�#�����j�����+��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<��Q>�����S����p�m�("�n��=Rd�,�@��e�3���=���|�~�[�L-#9�E��C��c��*=���M��G�����k��87E*��*i�.���VN=���0HL�A��S	e+T�=�*55+7��gj�dX#D�V+?�_L� 9J>Ϸ�~>eTt���y6���~%1�G.q�g�m��oe�RT<O��>�NV��RR��6u'��}<��o�0��H����	Q0����M_��at��н_b�""v���%'���j��X�ĢHI�'W̘��u�DOų��l ��Q�/1<�%�3V����GY��P:b3T��W�}��� ��:,-�Ϣ�523��1�!?ĨK6�D�M��7AP�Z�b@C>��6M
�;knl5-����;OF���D�p�B <��D�����I=�*�� �����!�~>�֙��½ՈU;��XO��hIu9߷qBp�S��J�%�n��lqg zE\����1� ���3����.|TYV)A���2���k��&�cZ3U4��>i��rdr|���B{i!�� �A�//oC��=*T8��]��eA>��})�ĤR��U�W}��!Q::lK�n�qQRQZzq��GJ> I�	Y���H���n\�$��̿�����2'G*�9 W��;�K��d����%@-~58n�~
%��+�(f�,�^2`�W��{��/�0�RZ_H��?ݏ�~���|���p�qͥz�����l�I�l\��&�*�8���qr�I��6�c9?��z>�>�2�?�:���ۆ{ C�1Ċ���zS��%}��&��p�ڬMaP������u�$��/��E����t� l�'�C]���ZV��< fj���-��S�>Db+�j�P]V�n���^ ��j�O<nYԩ	���+%����cǽa�EJ�S'�7�\L���]"�A�������_ؚı_���}��W����Ás�ƿ���47-���̽��H���u�h-<��ھ�JI�B�"Hg��#I��g"��7U�-�B/A���Vba\\|�h�H^n����1q ���$�ǹ�������V��lu5�t�uɆ���v��	�{P���\�o{�e����c(��)qAF~����2�/D��(�zq4ys��]ӶA�O�eN,|��d%�+ȃA��׺¨B<+ϫU�M`�փZ~��Êo�GcLih���gf䯺�-��vKvY�q��*	����k�pCM�f\Y���D�LFu�7���Jk��W�%�z�M�]sTlNf��@ ��`qk�->
����IjM�8Y\� >O��i����"���.��3<ᗒ��)�g����u���c�]�f䫸>���+r���g�cL��K��qgLtq��b�{��p��s˂"�O�;y[�F���g�օJ:�X.-Y�k]hm�|��azj��)D!�"V����+�a
��+1-�Q	�ְ�B$0h�i�y��}DAٙfue�J�c�0����!3���m���]�=>�� }�u�x�\�G����� ��S3�6$���_�\L�}�;�k[�h�~��A��B�C�7v@�<R_��ü�y��׈�_2���8�i��Tj���W\�h��*WRQhEzC'���}�?�{8��qkTa����v1��F�� �����$�<��-�������XFv2�-Ml��Y݀��K닏GG��vk�`/$8n*���n��5�I���?���=�Ϻ��{lO�ߒ�a#��"����[��}o�Y�?�������0�0fX6�w���z+�Zl�k�"%緓h%O��S�]=�g�G�B.8,}�������K1!T*6�Dk����R�J���:�1i�6��˽,^!e��[]	�z��Z����6��ξ�[8�ms��A���Ь+@~���I����P���o�x�,�ۯUz���gcjJ�U��n�[�����-Nt7:�޻�'����Q����@�����r�.����z���V6"l�����pB�e{Hi���nÁ�W�c�*.�EJ��"G���V�H��v�Q��áҫ��"1��`���"�m.��,	�.ރrg�/_�j&��vlv�<�5���Aٲ�}���g���2�SBg�kA�Si��K���@��b�C8ޡ²�D��S�2��?���3�>(tl�i�v�D$=���,��H��D���ݯ{q6��,VЮ�oĆu�&y0�QG�'w2Y��7�g���L�����xx�`Z0��
��}&�;[�Ѣu�}��4�"	Lht֟�T�[�VS_�gj.oK1��<^zz��F�K3-���]�w\2�kD~-*t� ےN$(���h
p��9�ߓ@T�Im���X��jo D���i�E�Ukd"m�sܗ%�d_)�O[x��+����_���?R��M��O�FQD���<�����LJ����%g���ҎR�n�Ú4u&����Z�����+� ���u��Ǟ&OD�-����:��:N��E�<��rιs�m����n���=u���-:���cmU#���90�^���AMM���� V���W�x�%։��ҭ�7�K���` ���]>���q����M��Ǝ�n0��D<�7��FB#�-�[Xؙ�=����
7��:aZoa�R�t⧞M�����x��l?� ��.5�Ғ��0ѳİJ�#���^aJr��Z���`�����iqZ��7	hnd��D�T�qq�|�d����uma�V�L	U����������&�y��A�V6��o"ZA$)(Q9��'y~�ɣ�5���S}���ZK��0��g��rƻױ#i>n�C������@�m`���؈�����.i�7�g����pK�"p���1_�vxo��r��a�g�|�*μ[���)�b��Pk�Ϟj�)�?��D�C�}��BҳFOà;�RJ�%�i5�Z9ZQ�cg'�[Y
U�O�fE`7�bWn�u{���M�\ʡ^��YH=�����	G-�Ʌ�����f���
/;����ޔA����&+�:�:���נI$�N���q�\��C0@�7�-h �]EE F��J-,ad�b9R�>쮆�}��YN�ۅ�Nr����5T�P\��aȩ��yH��.m�ʩ�,͊��h��T�'�@����ȶQ�Ҕ�����J�s?4��:�I�}Sv���G~�*��:K��Ɠn�h��݃�hy��[e���E}���ů��C�����s�]���pa��J�Ӧ7��i�C�,h���3e�w��y��oU�I�U;+�% �9�W�5+�8-em���^cH�nI�*�^ �țS��n�_�[{h��I?O�3lomD�bw��5(T�l����E���{���1|�_y��ܯb�1��RLPHh��h��O��	�A�dHo�:�7���,X����?��I�%����)��ѹ�S��9/�V+�w��sL���Ftܸ�A�_kn~_�+~{�,��!�	��`#�P�qk6 �;�2�����d��f���F�Q�̗�����16x��g��m��:�MG+��2�I<n͹?���\���H�'��92u����qB���uq������k&��l�s��B�;#F�}\gD,�hR+�@MF���p;����.Q$;�	�+R��N-HG�Ϝ؜��sc(����*$��l	�E��=��X�����8������%0C�T��i]/� b����;Ԏn��ٮ�8��mnc�̮�> ��crW4�*u��� Y������a�Þ�+�l'@`s=�����!h²�+���=F����FLT��3�sSJ���Ѷm���y���Bϻ<>���$��F��l�O�p�}&_#��q�i��_�����0�b�.�3d{��>^k�J�&�͖��}��}�8�8_�k)׌nH�ۮ:.��V���3�&qQYg?s�-$l���>L�|5踆�>��/56�|��Q�9C�L��-Lş�>�5�[�.:���cUt˜[y��W��Tƕ|�!���0V���?��4W>�i�F��'焮���-in��TKp������{x8���=��
5������ē�	�[��� Ľ��Q~9���"���t�M�����)b���c��x��p��@��p)8sX��%� �ju1aHܬU�7U���8��9���o�c��l$?E][4�|��KU����Ǘ��+ҘA���j�0��͖�$�F�[?N���g�t�j%ޮ_P�	g��u�*�Tk˯��%���)��)�;���?^��L�����BFF�ߔ>s%0{떰�L}PzQ��D�U���~��҂�o28�|�_C�hͲ�� V&�R{�ʄ�w�< \�0��	T���A��7&C(�7Ҽ&��G�N��]@yȺ�7���R�d�ٜt@�{0�tz�f�]G}J��d(o�
~���Q����Ʊ��J�]��$�j,/g�0��(b��OjH���-��¡��=r�TR��J�
�j����L,7	�仮̳-|.Ӄ���3�b�]�/�A�[F{ѩڦ2n�-���T*�v�k,���/PBE�n
P���h7i��*�t��I nF�\�R��ʈ�i���w�7$�,G�o����<k�-XS�M-@ч�ђ��[�މȣ�>�cw�ىöֺ�˘�|���W��Ř��Ч�[�񘵂&Af(�`�ٔ5�8<W�~/�����Niٿ�8��|H�Y&;�u���I�_NR�j' (��K� ���@2�)�=X�;6�,���ػ>�{W�\
�]��떂��y!��:�gF�σH��Bg>P���~{�`:0��:����i�Csk��p��}t@�=�S�&P�䔹�Q;�g~�߰���@ G�є�{����Z]	T��������|�<*�Oh-l(
a@f�g�3٠�H�E�xrlE�.��
i�K����Xim���i6��bM9��N)�w�&�%E�֦�����Y�8�i��K3{�5^�b��%lY�����;B@��Z��1ͪ�v!K��ݶ�+�*�`�X�0�u~�'����D��Ly��`�TS��.SC���k�����5�ilUT�/�D�ĉPW�@ȅ`�Z��ӟk�ی�"$�a�1 �\���Ů�,~:m�Y�fQ$:�'c�����!.+���'sG�گ)\������c�J
�L�Z� �!2_Ē|Bx�1��J��v<
E+�k�8�ܼńYC�>�=A�ĩ�%�Sn2������
����2KI����'g�M�oK7O�}�)M���bF3� ~%u����KQy���h�;�?���}Y�9A;��+��b;h�`��c�Hىq�n�QaژP��t����А1��F���wH�1!w֙4���،�&�a��_Գ�59GkI�/|4��'+v>�ڊXOBh���C1N�"��X�"q6ޅ����\�Ў �*Aۗ��s����
����ɦtNi����<�[� M��N�=[{����Խ�=;�(B����p��Hyi�`~<� ��mr�tT9��4Cqآ�oC�\��|X|p�i�<bJA]�]~�����3���(����p/U=��K��O�Vϴ��������F6�ԭ=��9�6k>,Q�����H!}��ER,f�|.�9'=.��-3��o	B �nt$f�A"��(5��q��p�~�+Y���s�Wn���J(���L���u�mg4}Jk� b���E�, H��M���f��O��Óۏ�le0���̶o�s����`u^��^Ԛg)C���7��*c�$���G�'��r��~ά.ń�@���hAZ�k�h�����<|��7�����n�E���a�(�m*��6-r�'�Of���Q���]I_�(S�a��I?8%q��2��x.@l�W�RO\��Ľ�^,�p�/�e�����J0S%&Tvs)��С��_"Z���7ō��l���2I<���~�Sj,������u7��f�c���P��%E�vEYU����C٢����l��1���u���7���Y����&[Z��A�%�+�&���^��4���&�PK1B�݇��m�$_��9&���&�ቔ(�Ƈ3����C��9��
`����A�*�n�#�����E�$I�^�o���k�F��O�o̾��ˀ&�����>���Y���j#��R�R��F����?Ol`�*Ǭ��������v�,������N�� &1�u�%�a���	]�̚�Y��2�`�޳���<Ga�͌@Y����V�F�ne
�;΀�渃J���*]j�!� ,D�����A�D��)M��ܖ�%d�_��8�H�i��P�.��X��R������W�9���c�큐qX�D#�%;Ou���?��/%����T�uI�btҥ�s��]�ߑ��ɽjQb6K|F��'� P�.pJAo˰]�ML�ZcE�a�P���9W8�'����4���ή��X�3�1����2�,�v��*��ͦ ��i�`/���rf4��g�{T��F4A*d�4�x��q��+ x�y L[��s����#ͤ^���|�"Um�hu�SL4o��"�w�i��bI^�GEv ��rN��"�v,.�1����2ם�'����6�D��<���a�>�꿨�M:�3(:�&}S����$3sߍ-�R��`��y�x��'�� �j������N�pN�?T� ���-�y����Q{���ٖ�oaC঎)���PB�@��h��8����QS�p%���;;YX��ڣ{�,��P��?WM���Ƞ��d*\������S�"��^���S���Y��.��-�Br��j;�ψ�ޞw!㋽�d���\�ݦ���e�;�$Lʢ���m&[IaP�g�׌��:�����О�#agb�J���*���`�XM�򂷘m����ǽ�cYN�SŗטAZ 2	X��w��9�_ww*����'���W���"��Qdh�0
�q�%~��+G�b -�������?;g'�W��l�'Ĺ�e�*0Xhc��x�����'E�x�,��@TQ�q�B��f���Α���ٹ����;&��!uFL��g�&i� F���Y_�m�^t��>(*L�x�f�'�I����%{FM�#בI�~s�gF����[[I]y���-(�E
�!��_݇(��zA�
��b��C�Y[���lwu
W���⋧�dbķb5N8������D�(�������R^U�Z�!'F�yN2���f��Y���UQ��cl���� �Pjv��Bʔ�ˌ�����9�F?ݘ�#�`�t�,��8o��l��8��J�ަ�1[���Tyc�\�9f`��$E�L�:���0{�������bfx�'!E���H�����l;u�ʙS`q��ҜU[C��72Ù�[��Kᛷ�;X3b�'+�r�/P�k�2au�J���6K���aӾ�a�ţ� �M��P�3q�R���Ru?��m����>I��N����aU£�)1�n�_x �g��iĎ=����`5zj�~Qq�	����~����ڿ��&���T��DA�!�_: �HT�a���O- �� )�/�b���L�(8.6��r*�@蹣^�ж5�Q��i������w������9�կͻ������;Xį������� z�
��#��Cw�^_���N�GzYb:�淝�ޥBBK��/{���u90���I�҇�w�]����"xC=���h�`�k�$�5K��e��V������+#	���mY��!t��ē�T��rG��1�5�aG�=�&́��lh63xc���E�\�ʟSŞ.��o� ��������ẚ��n��П�_�dCr���mu��/mq��G�����=Q�B\��RJ9WE>:Z�!��a,�bm
�dh9:b���D�MH�]����,s;��IB�r����ѥ��E:�sq�2��*�h�LM�(��`�]ig�b5�p�W_4a+�g*���a+U9~��t�z<�_�P�̩��P�B����n�0<�<�1�?b��1g�b�� �ۄm��x��vPi�5������Ԧ���nz>�7�,or�Bb��/饁�J���.����/0=x�;_~�kw߄����6/�hU���DK3��>bC�`��&��\�<��C�@`�/CK�<���߱xY|��l�\H���o�8�ټ�#��!�//+�
d�6�e����]��Q���많���H(4�Zd��r�8šAA7��(�!esը{?��蒊l�S�A��E_}�V����Š��17���������z]�皬M�NQ�B ������Ȍ��������ٝ�TY�%�����);��F����p)�^�P�K�Y��Rܗ���k����x����W���+j3�vD.�^�ɆT�M^b'�HN���_��C�h��	���0��S����%Z�S�u���j���T(�nj�mSSK�8�q�f�;/m�Ac����i�*�B�̗�1%�pET�6���l�v��ɢ�� ���d�y�;s�
�"we&��L���(��tb|b���ӷJb.�a��<�����`s�u��x�����/�'�������ä�	l�Jj�ݖ�U]�I�Kt�����s2b�o�*�*�2
j�C�B5eg9\0�}{���`,�)}�\p����f:���E�m�A3�㍛g����,(�Q/��#�Q��������ju7U1��2�rH$�;��K<>_�vb�X��ܯ{0�>E)���d=� ��Q�}��&MR����U&Q<<�@e���ʮ*���� �>�g��Ӷ�h��>�ǣ�JP���K��Kaa矽�u�C�T���x���Ґ�f�B2���
RGq���u�h����P�����gL�g��a�y�Y$G�Ll��ļ0�(�a��#`V��Ȅ�x�D��i��mG xϵI�O�m-3�\jo4�mu �7�Or��<O���E<�i����4����)�U^rxBnX�&��Y��Bv�{���S�μ{����%V�Yh��:�NJ�!}L
���g�����A� �2Q}3=@�mר!?NN����A��\3����ܣ��ƍ�Tg�
)G�Z��p��
K�L�^xe/@:�8�K��%��9]E6�hZ�'%dFѶ<�s~��<F����+>y,khH7P �8H�e	[�^�'o�'��[��Ȅ� ¿��ϡ��Q�C�z�؂T��Imma��vD��g4�rMK�:Q���&��Ʉ���E=��)vg�B��ѝS�Zcʍ��k@��%��ni.W�\�t���!�)���w.�T��C'Ga��P����r�k�0qnHڔӦ(�q@	^�!D)	�P���<�E�B�[�_�]j��;�E�T���Zyb��`Yޑ���!s�������n�e��ׯj�*��?~�� ��4�*��:�Y#�#$��5U#����|Fu��	:U(�D�C��|"�xz�?�4�@PA��I��_��-J��{ge���jP5�lkԤ��4��'8���S�����r�C��d�k;��|�(D߰��P��͂�l�5G��R;¸ۀ;��`@|9��+���5ܐj�hFt\��}+*Xx���1UOkoB�&�!�j�-/έ�u��rj�W����T�Wm������H���N�jH1JT�kN+>�ٟ����dC#�h���K��Dя��F/��OKW�ku�$8�ֽA�͝��ƻO<K|��&}��;Nݐ��~��X�l���T��a�	�n���{��wΞ�w��%�0�[��k� ""�w����~q�HD���p���(����m�����v�/z�,���:��>o;wGQ��:��vN�����[����x^��V�5���ʍ�� �L��YK��nySՕ��FHj��P;�)�-�muh*�Ku�o�|����^�0��;�]ɠ�M3p�qR�ISu���K��~4��Mq�&�}I��P��[ ����{:ƿ���O�\��2�����dcR9�S��80R�Po�`Z�Ϊ6��e4��"�C%�ooPx����d9������؎������J%7��(p��2�m�Mv�$4e�!LTl�tkc��G���`[;��	Z1�n��hX���`��">�VqJ���Z�w��ЬZ�8�P�x����mOѣ��;��'�`�\����d?�c$������R�N�pg\�<��WM�g�]�4����=q���d@9��"-U?�25S��0�k,v���T��o3�@�)���JF�t�ޢ�Ȼq)���_7���tn�s�:
b�C�i	q�v�*gS�Z&�i�h��C�iwns�<�q%��Ag�)���J[�S��v`��E���Y))�ԓA�]	jǘV�F���HM�E<������ТA�f�ํX|M^����#֏	A�����P��mF��79v9'���*�Ϯ��&\��֍�U
%�Q`�9�DH�Kݭ�vq�D�X�	^�HYd�kycwY��z	.�*���<���Yb9	��N�#���k����<~�\$�'���L��R78�;��6o��o����t�Y	*ݧ�a|h�b  �l���67ژ
�?�/O�o�מF`>�3L�^�H��ƨ46{_+*m��4UxV��T�������0�V)y��^��V��P�ӈ(s�ߎ����^o�$!���Uc∝����5.����t����[Lh"I?ܤmM�
f���#'KIC�q��U�33�C;;�뾡u3���'�Rr��������Ճ��������>��$�8`7���/�qI~�]��$��0�(�fv#����#��?J~�١�
��﹑*��O���@����i��b�@iw
Z�]6�AXQL� ��h�C��Xěl
?���a>��C-aj��J��j� /������. �x��xL\Q-�-����T�hR�q	Kѿ���z�-����p1+<�0� q�1�+ H�d�rW�VHeA�V=��?��������.iئFUοTnaםo-�s���>M����O��������,�M�N�=�:R���^���Ti��2���l���e��aݕd�ZAU+Y�T��,�D�����h�)��a�I�Pϼ�ɴ��c ���}�;h�N�d@<*��σ�V.	���JXo��q-��+�cX�!���^�|�p���8��[�4 j�K�R�{���()Zp��LGVT̟ԁN�/��?�Ȯu9
�(,z�*:Q�)��N���B�e`�jN��N�E\:����#˯����8���LeC�0�d��FR������}�@��/�X%�]��;�*t��Ԅwd:�[b��~F��l�\pl[��;���ٹfs����M�ߐ��!�3��" $ ��h������$��Z��W�&z��Ԃ��oH�sݮiђ"g�34'��:���3ss\kJ�Jd�ٍ���P�oR��ihIF�!c,��+&��Y.���S���UK��}����4��9y�;pbwtj��2��u�W��vf��Q��s���Q��|*s}{�X��]�����[�7E��s�{��s� ��,�L^lh����;�"�9	�w'�s5��O-t��7��~�]}D��b"�, ��:���[���ؔ��M�Ib�4FCF������5��F���>4U���)�(�C.�����A/LRB_"�"�	tp�F%}���LV��Px?#��/<��2�$8!J�h��"�����H�s�Ze��$m��� n��$�5]�)�>��Y0ސ˵ƦG��yp�%BMS�A0�S@�4��l�����{З�ǥ5�B��}�x�W$"�u�8��8��b*���O���0���5X���?_k��ь{��~�L2:�	B\��^�y���}]�h�#)܆vN��z�B�5�6�i�؆Fx���p��c����S�D���� ae���g�H�e?����7@	!1-�Jw��A�~(�P��p���g�?ih~��VZ\f��ܪ�ࣖϭK����s�܇ ����fS������l�4����A�� ���}7���1Y]λ�J�t����rG%�-��������$@��	��yG�)T���ڬ��ꖿ�RA�4���^�!8���zJi��Nk�4�_d^����t�F<hy��84��F.�V=��u���cU����̡,Xf���L������#C�a���Ё�_�f���5j�z��p)�]��VK/]q��n"���Ӌ���_ڢ�έ���/��R4x����g��{��9U~�0����6��.5�aK�V6Fh�e
��Ae�<��O��l���j�G��������"�Q[�ǔg�19�쎌'7���F!�h��\�Q�Z�M����,2;�3�8Ȕ�c�=;�,����|��_�HIh�Vt�zs���O0Д�&�ҹ�T5I/]�}?��~|Y8z�=/WC܊��s���3�'��l��8��e�C�Cׅ��Ds�+��Cͳ%	��k�����T)�0T�1lv`��',��"pw_s�Gk��9,�$��w�@��{�����&�6G��Al�43��-Xvr6��tOu�d�V��k����������iT�����,(��^)q6�|�WGS�ުH�C��;b�r��d�芖�~{L��2˰�E� �����YN�גM�|����Dkx�\�f:c�?7U� �.4�P��u�m�rrɳa��TW8�{l立����M
���]bc�9OP�eP���ݮ�p�m�V���K�:x�uGf�A��'��X^'Yqジ���8�$|�s�;F���J�dK��D��Kj޴H�G�[ԯ��6��R�,J���$���qN�Z r%�s�n]˵��@��f(�v$�ʒ#�M���P�=@B�#��6g��Rl�:��"Dx�>>�f��FaxU^a� �kH��t�|>n�PE�LW��#�P�r�}�?�6ʙ5H8[�!4p��
@W�(zo�raYS	erx�Р����V�)(�]�����jE/�/^�{	^J"rL��ȡ󰲯�Lj.���ޘM~�4�	I����)VU�g�D0M�X�40�hb��P���d��Ķ�Z,���K{�6�
n�D�#CT�DD�w���e����j�w��� �N[���:�Y�y�`$M2m�"��7��:���SGt勖S̠��J��*�"� c_J���֙P���o����W�M�+k���"yi1��}�K�0�+��~'�쫞ݪ�C�%.��6�G�{;�p��BA+_���
=eLgc���=��٤��\�R�m41���	��$�q�b�7s�\��g�����H�i�k���|��8���o��]�QTV�y I9W����[9Jk����mFBeB�l�4�&E���ږ��@R�5A�Oz@��9BkɁ�;�T�6�d��=��b��~�˼X�ٽ��D,�ƕ����i�<�@�#�5��J��3	�|�mp2�m�-ƒ�RQ'4D���c4$J7�O���9'H��)u��'*�����X8}�.*�|r���v�*�Qʮ �����|b�(��G�ޑS��<�n5_X��B�A��[��dq��8,�M�����Wd��6!���a�b���,�E*xIۉb���~X��ŵ"@K��Y�z��{Ŵ����X�T.�́���t"5(�2%�����<� �G���G)�E��������� h¤y�#���-oo��֑ԓ!�i�>���S3\�jڹ�._�ɮ�n\���f��Ё��BۚXkK��]d)%&'�^��*�7�>�י���4����l,���?PV�󐆦�>��(�=(�GȽ$hu~`�+ĩ��}8���B*�$�k�pd�8цl2d?�#���8�6[ƿ�)�(���:-��$)���C�خhSb?�E�����NX�f�x0:�z��+  ����!���rzؖS��V��)�.nV�m�������u���9�]&K�̳���`�ư��3�NT�w�5��80��3ǀ����DoGy���a^�p��(�(�g�\�����1>(��i%W�G!�mf��9���vb�z����/�<���m�,g��;����>��Y��$��m :>�Y��QD�PJA�S���;[�D�?��g�t��*'�iT�h
�`&� A9�C���T����SǤ&�\f�[#����7�w�^���Xk[|�9����+����q�Nr�-��Q9H��p���뻆�́�	����,0IZBCץqW�٣{!����M+��B��m���3!���Dy��CoTҠ�H�yy�b Ξг�4��W^8�&�&�K[��Vc={Ak84Nq�������5>H�w��!�\���5��{b����ԢV�[)����O���ؑ��+�! W�:(Ӵ���J�*��ydxl�0�{e>�#��PkSy���Z���K�D�1T6��|Fv3��G�i��]d�W����*kf�g���B�|�/#❞풔�9�V�R��M:%��?�v@G��^��`�ePow�Y����{=OM�Ѯ�I�������l3�w :x���CD��t��F������8:jM��\Y���h�3�q��O�Z�m��uR�_�������f���.�5�P���3B	:�UV9^I�J��a�Vp�]9(�`dS����[DSJ��4=�\��M۷���8���������{�ް�h�78�>0�6��㦓��X�Rt���m�ZvO	�×�|����帺	`0fWs^F��bM^�"Ԃt��}�}�xk~� �}X��ݙ� Ӑ���Qa��滗��.�|`�X�zk�~Z��/� ��]�j�e��l�)+�MsJ�y�QU�V�VC�
ضVn��jv�m2{U������k������9���#�,������p�5	Fu��r���ӻ{�y�5�ͥ9�5g�HD`/�����xJ&|�}��-Hى��) �
�(34�����n���/?׵��U�M|�|>���sc8��]ZջԆU�ms'
X�=�Y�B���Q3e���q׮X=H�-�1�u{�FY��`��l�$�V��F�׭4X�zt��;��-�m`��QWt�x� 5_3z������p�(��*��+��"�y@W�3�9E���NӠnw}��զ��o~k��I|��'��`mWS8�#�h�77o6Jۅ2� �!����*UA1:P�+ͧ'3���wǘ`�Ϣ�.���,���}�5Z�?.�Č���%'#&(T؛U��ݓ�q��u[IL΂�Mlrی�����1NV㻼�.��M�y۳?��I�B�?6L@3�5�ª�i�β�<yka'�S�׻�l�{��H|h�`����ģ�+�'�#��$G���o���P�`��tt9�G3�)�3$�L;tx8��a��f�My��`O���󈳔N&V��qFh�\\[�(��z�tXto�*���rt���l�	-��t�!��`����G��=I4�X�dI�M��{_]�?�$��$S14VN��Go���w;��߹���q�q\tb5N�/�GP�M��P�m��D�G*x�̘[ҳ)��z������90�ۓ|ɞp���b~ٴ(,��y�޾�f���7w]�$Lb�[hK��+d-�,=�Ě��P+Y��$n�y.�9�QK_�7�<m����
�y[�դ�X[E�w�H�������%�<�G�O��!�J]�5��W���������5ۿ�"gL��� ��#Y��WҖw����̾|����it�J:�������M��\�Vz�'��F���[QǣԎA�j,ʟ��v�cB7�>� W�3��$%]�i��������4����|w�K�ho���P�k�b�Z>�m#�����&t��1�;#Eg��T^4��0Ǔ��N���s6� (g[��+*[}72�F���E�@#��t�HU�w��� ��v�`H�F*qv�͎|c���ϙ�on�X;���fu�)<"tj, �>
So���軨�
����Vc�d)aJ��2��������O:���m�f���p�e�d��G�i`�¬�˒�~�)���8헭2��|( ��KJw��Cc(B�Q�d����e(�v��sCLv�&��X���S+�-Gѣ�@�}�%(x.3���g���o���/Mv��:]'}�񮂟�X��W���3�Ço"t1%��:��_��ps^V@�!	��n>݈7�l[g�\VE�k@�h"�.��˖_Iw`����?�:�H��h��]^�M���� A0�\���.��p��5���4z(��܁!i ��+X�93\ {�S�Q`3,��a���{�p����L��С��0k���X�F#�x����|#��\�]��k�ճy��R���3Luoe>8��g�H.;�c۶%�`0?�@ �O�+�ve\���Գ�ճ��و��ѭAf�����>�w��ź�Xf�ڹ���&��2����.�^�$�cgAڱy��I{�r; ,�t�/O�x��Ov��u6�l,)���$f˞�R�6��N��mhO��Q|2_DJ�t�oy�ORX�_	�{�9�ͱ�������S2�"���N�AQA��ȱ1*O~�wW������;/��e��c�
����Z �ȝN{%���$t31�G}�|�0|�9M�-�<���2;�l)��s��ҁ�ZN�k-t��{ze�P0jthT��!�ѫK���3ގY��25��� ^D��Rv6}�-�_ޖW��"�Q���;sst�����(]a$�uQo?�BIT!9�	�>g0F�Fզr�b��r#J���$�����������X����H(�Aʛ��u4Y���d�eW�XF�H ��y�YXb�;���N���1S���= Us��E4��9z�,��:yaQ<���1t��:Tt\|Js�s@\gח<��iv=��~|!��9N}D	64� v���Z�p�]�E/�Q�s��2޹/��b��<BZ���Z������s�uJ{��cq�WC}
{%;W�H��ˋq��0�����W,N����������L�/#�OT��6��	�埋k�F<M�Ǝ�z��U�� �,:aom?΂B3������'*T�\�Ok�;$�Y��e�cU�{ب@��v=�H���Ȫߵ#�����WJq߁w2NFp�mC�j�N�,G�ȿA�J,�Ɨw�}����$9����j�ޞZ<j��!V̩��4�S$3�����)C�u^~���G�K����+�A�"��98��x��c��@׃�����E������F4E/vn�̈́��o��bM�$�#����s���������gqE�Q�2BOC�PXҒ����\��9��ʽ�М V?�v�+�"�L�����*,vqc�����'l�߆�{ͣ|,�E�DUNꦄN�G[j�&�Bv:Q��;�HrR�eț[�YUS��*̉�2M�<hDuE�_w�8���
X8v�S[�
8H桦�"f�qg�mEiĈ�u�k�*O��D���n�����jO2�5"SU��{N�TAgHy�/~S��M\L�{w���	*�Q�q�9�� �n��)�X�x#�L�
�m#O~���Ae	�20��@���H]��8��E5��?�r@I�!��!���fg�Ze�R�N����n�`F�n/S��E�l�Y�3쀮IY�m�� �۟����2����M�Jw��˫��$�d����p�Èf)J���ɿ����š8c�VS��i��]2,�(G���kJ/��p�t���U02�]�yM�,�WG(�<cC�>ty��� ~����lb�3R;β�'���Ɋ����l!���R���h��C��3�#��t��	�#���$H_�JP������̨�:�eC�|�< ����u޹)g(?Q�A;��H����n���%�`2@V�fn?�Xd|��'�7z�a4N��?��`�F��Zo|=�
��m�,ڐZ�l�� ]H7�_c�s�ܒI-YN�o�o�w�H�!��-+Z��>YW����R��Ѐ���us-��PH�\z	�#��O;��8w)q��\[-tJ��tx�o�h��%��Υ_��Sm/�@�e�7����� 8�c��Пm�MR���9��W� ���=�{����2��8���t`��ﳭ4S�F�-�
N�%!�j�}�ݳ�U�!�^1i5��SJ�K����l&���6��D���\"���3���!��{�蠶�O&>�X�W^�ˡ����^�6o'���/�t����Hz�;����( �m���e����s6�Ư,gP4��3v3��}�2��l�B�;���(|�t	��ye��"�6Yg��F�k�M��"Tt&����AJv#�/�UȞ��Z�4k�p�D�5<���K�G��@�9����Ƕ.-���L�-s�H�=�h�p�b7'XUC`��w�����h�4�����~E���R���6��`E�U��5Ti�+�*>�k!�?�l��ح��F<�p���SU����#���e:-��U�PƼ�"c�&�� jp�����;f�OB5'A����޶87>�V��>��|�m�-��e�ȿh�8�d�h����9ޞ����Q�k��g9���B��������O��.~%Jǋ��MbkǠK�+�K0(�%�C���*��ɑRץ��Q�5�]/�噾�`��Y
�v^>�U�M),͌��^75��Cna�Ue�Ƒ��W%����z]��P�^PkK�U�]�ЬꯝI���vc���K'�X}�}��Y�lvV����=+�^�_�@�
��j�2G�F�'hƸ<%�;�XH9��I��L�H|Y��ϲu�qdWa42�n��]{�Ĕ����-���4�3�K�����'�ΜI���l,#�ig5���p����l�-�2����P'O�
|M�Ks��l�0�zH�O���U��j1����9�ϓ��XZ�C^̈Q�kB,�2��r�˾m��YO8���c�3�{WA���}F\�ї�R�[fR�V�w��+3M��p-ͅ��׀�P(�����M���c+&�%���pb$B��/�73�]&L���vؖ�\S����߻<u}���nW�������qq=�i�$�xiQ���`�s� y6��¶a9�� 4AA���4&Hw4����W/��5P$����↎y�[��P�"Jx��V�cr:+���?Χ7o91oR�X�2#��ȍ�V�����'���� �NyJ״E�{����	��_85ҙ����E�9��{�:�ľET�uA�������	,��)��*��2���	-���Uޥ�V����d�h�	�<���]�:�s�R��\eT��'f�Zikt�!�x����i�̗�5s�c���<�?���	\�����z�����8���u&�ĨsQ��M���<�)@=*7�R-�Q�����<�����Vɶ���ZG��ý���nB�ǌ�R�����M }/�;�n#�#�����M���׽S:)��Ǥj��b:2"���J~��m�]l=�j�Y��^���IK���MT��>�%�$?��1�t;� n�>�V�Av�۝"�ky,
�Y�:M���]��8�e�f�UR��Z�qt:�E�Z�G^*�/"G�����xSIT�J�t��4vxANw����$慿#3�m��*ط`;�D��(�"U�s�E�e�Ugȏ�y�2�u*=�ti_��JK�@�Y�{���B�}J��x�3	k��_��X���߄�2P�Į��/�E����c�9��5!�S`n%��g�v�$�r��5��u��q������q�:����c�&˦{����\�=�!����KE�2��dj@C��<��z��%��M����ay1��5���H!fS��~'��9Г���'��yX�b
��1H@��j���+��>;��fP(�IOEH�%�o1�;���c�ě�p����^�V�N��ia@7�Y�������:(Kҡ��t?r�
*BE�PgW�ގ<����j�C �U���Y�Ԕ�Ν�efh}39�%�j�(�yVY����q��A���n��	����$j�(%���)��ʹ��-n��Cw[�Ӎ
F� ;��C5b��P���g��Jߗ���!�ֻ�� ��Z�mbZM�2�a�4I y�{o�|�O����`�p	Ã`��Df�~D�<i�m�|c��4xdb&��m��IVA�v�&#廷��p}��_7�u��\�%&���?^��	b�Y��sMW�_Q����d���i@57bZU��]	�'�ư�N�]�q!A��_M������p'K��Sщ%�k�*��1�y�4B�������į�zʂ�	�)��N�︯1�O�MX�tM�%[��3tZ��[�Qa�t�{��v�ԝF��+_���g3:p`$d6R�	��%w�I���T��P��K�LtKG=��F�˳{t����Ka����C�k�K錭j�K~
V�o�^N:"U��>2@��/���:��u%��l���S�ð{n�����*��L�Q9�lU(��!���a�������M+X[�A���,'j(K����D@1iГ �a�Y,�P�w���2f+�=OC�a0yn�1w!�����Vm�7��������h���3.L�+��q�}=<�I��C��3��m3�r�c֖���`���%yZ��gT�E&l-I��yY��Px/%=�v�6 |��1%L�A8Ew�|f��k�����Ŏ��ϸ�Z=�z�9{�*77�{1y��y���	����NF����wH��7:~d�����qz+��Ċ_�����B�&߮C�A��ڶ�A��Z�E�#|�\�{�6��4��D��I(]b�ZHIX����dR�<�3�ϵ�[ Zvj8;�#B��� ���qC��V�KId_ww�ąn�6f�#N2��^-�L(�"=�a���>PD�(Y-gc\�ק��R 3Q +̲3�A��>�o��-禞O7RU�Ї�] ub�1�㊏�ـi�Mp{W���� -6�U��`� u?���V�t��tQ]i��J�y[�U�y��u9l�(��`�	������g�^e$�WKy&~��"�m��ْ�9�@�C��R���B��QۖFl�Yp��;~l�{�&`���$,=���d����I���	������\6�`�o������=���q�o�T�+h�U���=cc�[�s��v�3H��?�6�P�Ӫ@,��[Y~3(]i$����5��$ ˮ�����{�.�*^m���5�)��������~眘�m�(
���y��e{<Ut�t�T��j��BUP7����?ύ@H�}ŗÜ�ǵ Wgk?U�N����I��N�$�M�ު$R:N���Yp�Y�(o���nJޚ������J��n�a�O�����x��r) @�4
����EF�����1� �D:��j�JFc���R�Yᐿ�4�Q�B`�w��)��먯���m�$�n(z���C6)Aۆ`%�7Wi�!�AJ����Sw��no�W��&N���cr��r�ڂ�!��-r�"T	�M��q(ho��V��c+�Y���Z� l1kv@�|�(t�~�ڏ�����Z��v��'��|HT�[2�mD0=���@��-��te���\'�
=f1Ԗ��ZP�||p*�����qaԛ+q��/��%y���V�̃*QJ歴Vo1�5zN3z���f�Vcv�w�=�J�ݔ���ـ���h{�/|�+�_I~_��[ʸ�A��X��k=NBZ��2
_H����7#b-E�P�:��|T������;a�_�:�M��y�B*�[q�Ix +�o~�nX'���3���t��t�DH���B\���<
�L��x4���;�zL�Om�-QWe�z��UY�[��J��`����?(лD�8�gB����P8B�e_#^��h�cL�yk�p�(�D�&�d�'�5/4�Q$�r)�i�&�|
�O�i��R�,�j^o��d7iݽ�	�k�ߤ5�4��z����N�BVú�k ޏb��Vuբw���מ!Q0�΁�6�d�x\�.e�"��x�h|�Pf��f]�)�*9ʴ�������e�;jH�@��fu�74�ő�F~�2V�i	���so��չL���a���smd�i)�pݰ���ɽ�|�|�˺�a5�2�V8f�6��U � 3|�7�f;C�>8p�kb��.:�����I���NŀLs���:R�ͩ�k��9����"�D�X��������ë����
}��A�7s�S���� !��@�}�����U	FKq��G�߉j��!�T��V��+ѻ�=%�o�˧2E�etЮ���Β��_(�o
��:d^�F��۠
�=���,�m�J@8�\(��h��"��Qt�6	&s��D3�TD[�MK�Lɖ+�X�Ƥ����Q�<ը��m
�n)b���
��e$��r���r�v%���K2
V�4��_��}b䔡'-��
����o{�c�k�l�OG�L�MS@(i��idouL�z�|�W;.�[�t㱏���ڧ<H9$k~��~� rZ�A�Sc��@� ���/��X7��0�}E�=��H]���&7�\��8ɻ�-d��Ժd�2���SM�4 ��EY< ���EU�+�I�O��RtTDu��p�Jrah=�UCRڅ+���/G`��
��\�'Vh�0BZy�ޜP<��㷛�~�����%ȱC"8�}׈Q��V
�P y�<�!}��Y#�%��5e�Y#[���m��%���h�j�X �)л �n\N��x����:s���^m(k�����Ӂ8q�]�B�6��'�/\�zMɢnI��=� ȓ�g�<[���[��*]\�H�D݊���X��r�iȰ�|RJ�E�4����[`��S��
��r��	�F��#��݄bc�V����;��'ne_��DN�5�q,������$�e�"t��1���ɏb����:q��B"�RJ9}�ŗ�dؖ|��R�ؑҜb�^J�R��.�\����Ae�FU���7���}��q�)(��'��R�y���^����m�3(���KJ`R��P�=:���3v��fD�Mz�m���#�5(�r���h+'W���?tg/�/j�p�x<0�VF��S*��鰤���1�# [�vtI/���3�\e��"<�$y�E��|C�i��{C=�m&v	?��C3Bӽ_9��[aV����Go�w}9YFp��
 �*)-��:稳����'�����Bt܎�C+޹t!���?Vl҅w�8�.�7}�3LՈǔ���r8_��t���ܾەC��[���&��2���Nd�x}k�O��;���w8��m��!^��/js��
���ɹ	kۑ��J�?�����%��j�����N㣢�?0���{if��-^����(��7�����8`o�VeK�_���
��%��2���'���Fk�k� ���q�P|�Àq�^�x��g�eĤK�Ό��Q<�.?:J�ө���6g�=��)�zӅ��ųᬵ��}g]<��B�=���VG���$����3���#��b�_|	��ں)·��A�:��� �@��GG��(�F�/���	@�X5�]!���q��J�o��,��Ja�F��w����d���Ȩ,����X#A�x���BŃ��R�+���Fv�;��%�Sص�RUر�y:I��8[*t��z&hb����a�O�ڂ�-���u1�}��h/�w��~JsG�]<ǘ��77���2y�z0H8�H��+��"P�fpwc����惻�#o{���]b�MV@"��08"�!���ў�c�3R���~9Ec�Ҽ�v;)�&5�o�r��>������#���P��[���O����D�{����,��Jr8��I	��v!�,P�'�.�u�݁�rߪԭ�>,�ó��t�����S~��n�c���.�՞Ƃ4�%Ũ!<w�
+fH�����}]k�)~�yO�!'.5|����Y#��No��ƷHv�`ud2���J��uI�z���E�)[�&\���}�$D�C}�)�w架w����N����Q�r�:'r�FwXy�k�Cnk�'J����}��Mv�B�MAs� b�L�\I�jz�Շ2 ���P���Z�����q��h�V�Kh	�O�����eF�ޗu�}(SA�5�y��(i�d*L�3VB��?�����<n���U��䒨�h|Х�s4  ����7�k�8Df�D�P�q���
5193ٵ����#���i��PO`�1k.���F �̧�2U+�EM$W+:y����F��S�Z��ߐb�ձr�r/m&�-�A�����M��2��t�'WOV]�&���M��ǅ����ԡ(�n�����r�<mbʥ��`�O�Na�M� ���8u���,Թ�"A�IE�I����Q�vN��\_�������Š^;���@$}<42SZ-��.��ȉ������le�m;����:�pcX���V��g_��ػ�I>��%����(�{4$T �]O�N�
nmG�-
���#�$
��>�� ��΋�!����uVs���Ѩ�05�-/�)nth�8l�����	6{���<�B[ޏ̽��������N�CΖ�2����E[����ؼٞ�^��ӂK;�vԹ����	h��0\���v�B_���2b�pO���!�������٠��{�8T<��JQV���z
����:�v�$�PD���|�|r�u�(ϗ����x5��ɲW�R�J%#`oс�^�y42K9E��<��ǆF�p��B���-���}�[z��R�k@������өƐ�b�_�Dŵ,1:<�T�����/�G�����F�eVJ"%~���-�H1O:�Hy|F��nu��1$Y�-�� ] F�6���x���$�/�c���}p����8E �]�z�A8�_tb�-ODT��E?�	��W!��x�����˾��b�����КrػO�R�c>r'A�=�td��I9D��:����-2?.V�lŊ����|�����>n>i�!�����*A���O�A���}����D?1��:�*]�x�Ĉ�>��i��?�����@\�f��ꏘ%�2�4F����1)��<v��,���,x8�*�v­��k���p�R�W��?�t�9��A�:�$l��z|�����!U���M�g!���L�&�Cjc��l���"%h�5��/Z1�.e#�M�D�%a�f�\�弡<��&؞0Od$�� 	��Ѕi�9U3:�7�BM�D�Jyu��ݾ�����������Z���]7��}��\�\�H��;B/.��K}C�8&����ܧ�%�W����KR�{�m���N%0� �D��F)0յ�氊�(.�����p��?H�=�n1�#j/]ٻ��a����	�Q_DlT��
�h���ς&y�\��$HGJ�Z��luT�IZ�Y`r�(=f?Cޭ���M1�?��c��>&u�	�Q,0�e��I�5���U{O��{��n}��9,�R�0v��ta�����q��ڢlL��������T�����_��#V2���Bݮ?Q���1eHm�<�vl�(G}��!ե�� �Ϲ��%μ�f��i�]5�����,��ʉg��p�0�����ܲ�SC{��� �/6i2���e�m��Q1	�r٩���vന�D�2УA���X�]��/
�DG��$������C��+��<�{Q:���~���'���[+Er�o�g��UaxUˏ�����ݔ1e�v�n9{�����4��襙h�1�M%="-._5�e���CIC�����g���z�/B����a��`f�¾ �֙\����4��g��&��:� �MSo�o���΅���4H�*�eP!4���Xu��#Ѓ3ˢ�Ao�ʿ�����V�Ϡ&}�ҬQ���T"�c�9�*J,
h���3��W]�1�3�?�k��4L )��q�R��e|tHU�zE;��Hq}�"<gS壝h��Rk�Z�!�c�?V�C;�����?F5/涉!j����?� �Y�S�{<�ٛ=�p���4�z�G4�cV~u(�) -���j8��0<�e���9H��"��R��VV%Oq=����<�"�)�ģ�)��ѐ��:�2�<�C��w�X.��'L�Ƴy�
@���1T����dX����㰃�]C�P��zc�R����aཟ�ș]ҳ�82ks�v��(dd��%�^��Z�̵�	W���j}n�u����_�-6���c%cܼ���;����QY����B�����NZK~/��4��I�ф�t���>n��#�rY�N����_�z+~��� 5��f��j�/z�L��&vz� &����)K����BwKC��+�P����$�!#s7paIx��]������BU����+��(F�m����x��\�8wm+�B���Ƽ��e�+��G�|����	�g���e�0� �YXU	�%���釅��﯂�R\�˼Ⱦ�Le�@�U��VT��z�J�Z�|��.Ƽ����Νh6� ��h����X��?���Y�����ժyC��:�������4�G�AQ��4�����Q��ő�ag}�S[�Z�����G�́LMy�sɛ��]���qko�F_�k:����Q���AJ@V
*�����34�gB����p�t�~ �R��a��bDA:�`��g
-u����H�N7��m��6�[y܄y
��G��1ga�Q��3�:�T�S9��v2::ߒ%��<�����l9el�7�� e�"5*D%PA��v��Z�=)}�N�cW�zS��_��_ѹx\I��de�O����k�K/����,T����|D�n��e��L��O�{����o|�2Z�7�)O)���U?���E�n=;ț=���|k��o��"�{&Sܻm�[��#����A�!]�@�k�e�¤�xH��5��-~��Q������ e�H6��< XÉ����������ʱ=H��;-$wv6�MpX2��œ6�`�%-�O�ZU��{�({�Q�����e��{�(�B��e>��gX�?	���@����A7/�A�V`��h�O�R���?a<w��Ro�D�0�!]�5�A/��=�Nn"Y��C���-^�<<�ejF=\�r���GE�s�gz/�4`1~$/u������u:"?�������n�
��`T����*]Mh�v����[e��&�N��e�EY,�;����aj.����N�f9�kH6%/&��>�5�"�5wzm%j<2=s7+vxDf�Ʈts�)��3�Y.TCr�������\��RY���+Qn;�� x��U��d�z�c@��
Q�+y�������F��$ҍ ��w����Z1*�@2i��t{h�Ӭ YM��X��Rq�}3&2�����R�3�.y	�Q��)g˕��í�pX��]x�#����؏���>��3�p��;���� �Ln���Ĝ��!�J�|<з2�k��.\0X�d��}��W4�7�x�*S�I-@[Kj)ՠ`���c������R8��r�4�x ������EK����i�ק&�xPR��>��pm���� ��b��tg�֬b�yb;��ٲE������	��]�^#؅�Y�WgYM�/Z�z�lv��w�z=I���z_�pc֋r�����(t} .�I]�/T��hD�[���4�����5���r����f����su�8û�J1��A�-�����6�P��j���@%�������E�#L�"U�R�,�|0tY^�8��V =��dC�4'����x��h+}����)?��U^|�O���:�y��כ:4�ޤL�2��&�#�Ł٭���8�2���h{ @�B	!��7C�����v��NH4d���O�@� bKI�-8P\�����g�~�yd���Y�0���g���k�6�G�G�P���jU�n�c�;��G���d��Tp\<h���7
PlK���L:]=���9S1`��{F+���ۦ;�:��"U
s1CT�J(H��=}:�̰/����;2~^]t�wMA�~�]c9�Yʺ��6�	d���!���sM��|1b�&��$�Un- �XMkL���)i��ݤ(OÓ��E}T�>_ު�����Mh)౯��3����������WiŪp�u�2�ڱDj5� ��@�{��Fd��^c������G�� �s�W�AT��1���� �ړPe!� #g�I�,Z%j����m9��O�1B�9��)'�dq�6t�w��v�I�K�þ��N-�r����(|�=OO�pd\[A��`p�T���u�`R"OD���	f��i�p�ϕ`/�&E����i4�-��z�I�-ޥ䀬�GsYP/�JzѠ� �����-a���<�u��W˭a�����F� �k��8VX%��;��L�~J/}P���1xu��z�2e�9�TS>��9�3X��ρ��4��&�i�v��J3�el��p�V.�0��VY����$�%$24K�4�z��SSZ�#�N}��אRK> j+?����`�G��| ڠ|�B�>21�]u˪P�i�e௢���P�AWY��*���Z=�C�+�4w��Y�c,�U(�P.%>�&H��B,���,:֠q\�\_^�E<��e���ې�[z%/�3���9 H!<����*�����N��oÝ�b����02��cVi,Q��6�}q���Mi�,ʺ�[=]���ǈ~�.�G+[�Л��U����3.�,������~���i���HĔ��vf�\�-�EN����O'��t�Hu5�����|���'��e�Ok��_K����A.�}CT)�m��$��?��_���I�^Cg:^�.'G28�iNE�L#jA�FIE�/���8���y{�K���?*iJi;6�4��ǚ��Ϧc�/�w�/	O�8�O1�:o��z5���n���t����?'��M_��Q��I�E2���?!8m�i.�X�z	 �vn�����y���U.�J:�0�p�KA�X*�<q���z$�ۆ���Z��k'�,��(By�h���	�Od�zn<�)z���UB�G�Z������	��ͤ8�<�r�E���\B��ukxc&mGg�|)�>?����IX�V%��X;�ݛ'��X����S펙�� ���`Ԍ�@�$R9�wWD��Q\h�n:Kخu��{�`_~{�%aQ��`b+i�T��Ӷ�l��_�s)7.�n��d`}�(ȫ�%d������	a��V�����<���pX���oņeZ�Ѩ܅m��T~�$��e��ҷ������ �����3z�Ύ�ZW�O�bDO}`��@���3�j�Yw�P�b��ą�j�����2�$�ڕ�L�^�ȳ5�����)���F���4�t+p��P�KJp���|R/tt��=c'C�wh&���@�~m��ƭߡؓ9(�� >��}ҰF����^�>���O]�8,֙��])�KJVͿǖM[�T�j9�N���]aa�����{X��~�-.�mm�_�6nb�f�͆�����k��f�RPD(�[��Zː�X�(��C����a�*�t}�Y@�^�64��W]���f�s4��P��G)2!T�Y�j���ж*_�����!��;��8�I��k�=p�4bЌ|���Q�� kP�� ,�o���-�,$��,'�ˉ��e(\4U8Sfz�)�&k��͂����q!VV�잘De��@d���U`	n�U���n�b �<�l�=�U����7Z��f��Eʹ���7�E������� ��,�f[�bS@<�I�5�|�����Ń�J����q��L�
�k���jY7�Z.��PQ/��.�"B��hV[�Q)i�	�w�{N�n[]��(�ԥ:�%��׹ ��B���eJ��HD.�V/��}>hq�/{!��ǢqYy�|Y�Q�64 ��I�����1*�3���v�YB�;k����7�J$(Q�W�*��nLfa��dhJ嘧l3��q����`)o�����L�������	-�1q'e�x��H�Q�P���ӓ󨒥iђ�8�uxaZ1	8R�����.i�f�Y�ګ`���>щ�s�%�O��4u�{�y���H����3?�ZiA٤�#F�7{nb�\(��"�k�Dm�q��ӯ����30I�<�>�paH��ѭ9R�Ҥua�BRmT��9�n
5�n��Jߥ��y�=q �M�#���?q2U]��\u��$�NXq�����v�<�1��5h�Ț��W�
������:;��LQ������A\ռ/g���8�R)��Ve	���/�ae��M��8e\ ���cnx��^�R��W�!�騶`�BW���Z8����N�)�oaܜ�l�F̦�-��c��G%�U(*�"���>v��\�L�ƍ";s=`0uߨ��ˋ⵻�p�I����N��'�[��\�3v�_�����l�;]��
4˄,�[��^���W{���P�=7-	hU�ͫ���Z�(�c�L+���H,���x9��5�c�bc ��6��P�5�M���M����sVj#B�[�d����l	��&�	r
͖�c�sv���R�t������5�nna�M�l��(�s˽_�������6LTWH�� -�: �
]^��t�r�(:]�DMI��2��֢ �\����;�.�2]�����Gⳮ��qSE}��hn1�f��)����.�oԄ��3��t��گ�}�5�ؿz�U�F5D�"�զ`3n��j��B-w,�;�fC�c�Gt'|m�[90M�U3YS�"���S�QBӻ�刌���K(�݌�2��=���1�9JƮy�t�~}:W����{p�Yh��T�s�N<��G-�O'D�۩�
鲆�|s\�c^����u�LS�,A*�f2rʺ)gHVJ�Sn3��9���Q<����DA����G��&Ֆ?����[����c�Qz���x\6��}L�d���u:��O���dZ�EH� �LW����O,�!b���7�XpV����]|�+& ��m�KG��!P�����%���!u���L���֢��jA��&��E��F7�@)L6�4��=�0]��M0"d������n�r>�K�DE�˅��vSf-�S͒�ʽ����d>)���n<Ǖ�oi1C7
H2,�h��_��
�!:5}MOů�yCHn�i��M!�S����u�9�Bw*x%b5��3�?�ep(5��-�Bm'��h��ń�ik�>O�����YJm�Uq���������,L���A��M�O��O�*,�P�'����7�r<k�b��[c���Ԏ+H<sg�
t��AUsɚ�ƥ��F_Z���A)#n_����EB��+���$���䜆��F,
d�4B��8}u��\J�2�|�3�<��x�S͐�v��+C�Ky�J��g0w%����$Q�զ�B��!���i��4"�覂Lg�r�Z�� 3(-�Ex��"�
U`I��t���r�#�����;g�A�z<��]峽�0#L+��)��w����`$,�k= �T�w����]�?�/�}��?���	L�H���QiX�LIʡ�n����e���˔&������)^%eXH�#b�L�凶 �I�C�ޝI`hȭ�V���A2���N��%v픠��W���χ�ڣ��?�>�@�:�9��P�ݞ���G�M���i��0��%�1"��yEՋ�űI�Pl�K,HK1�7 �۵�aiC�$�#I��(>)Ib^���J�*�>���{��.;}�tޗ��r<k1�2(�D\���{�ߓ)GR�jVgYL2��� �E�~���*r�{{/K|PԊ��]��Y�wX{�ȗ@F�`�M�8u]�c��V���Mq=�}�r�g2�$�xt%�U�=����Z��z�=],K��dTz�8�����LORo������L�*����)����FH:M�o��A���2�­2�S��������L�b�-���[*w��U�3�r�pym�"�5�
���G�C>auHn��hi�I�Z�5ߒ�C�M�b���q� �d@x+�2 ��[��`�����+05E�;tOb2�h�Ą��VH�D�#��
�Or�S?��ΐj@sq�)����9�h�OT��·Y���֎u���S����aC	�%��֭!^?��w�1��ͪ��14	��p����z?�t�ƍ��_pa.]A� ����6K�ms}^��_JK���UQ�y�Y4�Z����ն�F4"me16y,����@r�rx q�.�oe�Z�h���+z������mT��@]W�4��P��TF��M6�o��f9��-�Z��؂���O_�>[T��@�Hk͑�A�K?��rS�5�S]�&��J� �z� �w�Rz�dt����_JPOD��̓�r���(�Ӷ;�!�!{�H�T$|�5�6��,:0�j �霸�AQ�3D������)�%����J������ \!}˱J�C_�2�1�i)p�;6Bz2���6�2ra�-)y�#�E��rIU/��3i��NP3H[X����b�?Kh\��p ��?�C��w�7{[�1N��E�!�e\-�a� g�($�l�)�����)�@�����cX��@�*�!@�-��F�ܑn������7:׳�&t$Ư����R��	�~2/t�S��8���sm�</�Yܼs�@�X�7੦��ԴJ�,(�ŗ/ى��\��BfJ��gkMu6k`��� ���k�^�9~9�~|����?5�'*�7-2+��A ^���ƻ��*��ON/��Ԙ�I�)�$�fv!'F�\;� �[�+��w����t�M������W/�d�o��\Z]�y&
7����c��,޿�nwol�6Fa��OvC�%m@o� ʯG�A��	X��"U:y7���ы�oI��~�o������d�n��{��;E�Ӈ�Z�1FD��7I�t�E��e��ؐ^��jk�7��e�Gǃ��P�,���"�&���
�tF�)�i�A崸M�3�_�AFh���n+Y�m���w%��l��q�!�h.�����`�ΛC(��B!  �RL�a�#i�m�m��`y��j"12����<��E�C/<������i�u�c����-sUI��1����t��(i��h���S�ƛtz'ߠ��Qs�k��W'��G��< �~�������|�UYV��d�����9w����'rQ��0���sc�^,��Qஂ����e/ky�n{��g�Q	|��7�=C+r��8��b���,U98f�w��ޢ� ^�'�Jl���l��br�k6��z�����>΄�1��ƺ/����,PN� ���ʳq'Z�P!!I@c�M������Aꀅ~7��Fω>�G^��O�ZͩH���y�a��O�EjfKս�r�xT��G�t��ΩӍY'	zr!R�P~)����N⦷���G8@��~���Z��% cN?�h�e���\)i��@����B��s����u�@�-��@I�eL#���C�L_+��Y�^�5E�1Q>a�m�("���PޓzY�������~�Z�khau��oC��e��s̾=�O��pSX'�s}���C�qqp�.�6�������W�];�I$��F�f*�6}� �ݴg_Ȟ��
ri_ ��O���ʨ����f�����!�����=�^�b(��<;�+��Q��3�ʯ�@ag{���r������ʟ@����pT}s��� �"���^}19�6j�i��9��Ԅ1�4PPnZfV��1zf�͋=��7O��ɸ�zX.�A�OW�dg����pYK�)�\Z}���RA˰��0Џ��t�YeV��ݔS骰8���Y��k�x=��]�]A+�02u���h��&�&�&�����ݤ�L���@5@cE��U?�D�T��(�0lg��� A{)\�=��<�sL!�5�^�B�m(
RM�	�+J�mnD�1~;��M�����&��n��([�P�Q`�Z �+��w�88猑#�Z);�v+��	}Tv�V�2�>����Ug����'VY���L��
 ���e�p�;ġ���"LE�۷TSI5SL��;O˺�??�p�6뷌���2>ۅ����t)Aŀ�ci,͌�tY�=2E"P�Ķ�ʭ��c���$�����c#�QB�+�Ǉ�����EЙ�Q�կ%@�$��Gp7 �꺡���{���4��zl1��	>]�8�q	�EW�����6����F��X�ea�+	�ᅔ.$b+H���-3U�s1���V�܉l��z����B̔�k"��ns�G���[u8�ku_����o�L(<�����p������epH�nnO�n��\\��6fJ�aP�R����`���oF�4n`+��~ �#4�-0�̷-�0)� x��f� /S�I� �c��X8��MS�]��^*�;�����҉e����Y��uY�<�q>�B}J-�h\�z������`*'�/9�C�3T~o������ ��6c�k�cj#��Qu?%���άx�N���"�N��i��(b���Q�}��ȤhI��_!m��7��D'{z�1������]Q�.��BЖ(:'IUj�X
Cۦ��XoHZ4�����%�1�6'�5 ȇ��K���E�
?d������
�٬j��?�a�lKQ�����:aUW�^SN9�c�m0����F9�nvNIB�䤄IY�q��*>��E�<x�I���W�ѐv�X����A176�|59g�o�S��M6��v��|1��8�;������
�W��ze�M�4��ނ1؏�W>������ �0����Ce��*��-R�}�g�FRi�d��	6�p���$ۖ�[W)�K}%+���v��ɇ�Ҷy����ܳ�E�Z=ֽ1J�1e�>uĶ��7'�\9�W_hb|�Rn(�M8����
����i�������q4�?�	�����{rP�����n@�������9_Ȉ9O!x���{ʍK���t�D�y�L���0�Zq�k�LMC�To�7h��ǁ�Y����=e�z��^4�/f2s� \]������XA�fV�9ꅛh�é���B�Q�2�Fnˡ���glY�l(=��A�<F��`�;/�����e��澀�s� ��ݛ�nS�"R��A�y&�Jk Q�Q:����řڥF3}B,+&�{�dT2�N�Sna�u��h�v¬w���y��\�^�T�71 ��)����ϋ�h��.s��Gk}�ք~l7q��HVL7[��/�R�X�v�s+�畭d����>ߗ]P5m���m�Y-!]�t���$�MJ��D4ݟW����f��'�j=S]��o�g��h�O����x��v�K�,�e������hr�❒�3���"`ygR�~�\7ל4 �2�1���x�2��".d�3{�����5���`y�t�l�H�����A�_f������eo
E���� %���I��4�<X�|`���ۃ`0JŮ��G}Q|����<�s��� ����S,��f���#x�q�����oUmU���� !���5�ߝh���O[�;����EC�ї�w$�C�*���E�{�,=�+���'$iN<��7��}sd�洡=�/�n�ķ,�����Wkm��c_A��1��kF��a�eg�'�V˺�d7 X�S�����������1��h8WkC�h�t�[)�F���"4�'�b�u���T+�|!@���wv���('�%ϡ�whi���_J �Z���ޚ�弰�nZCp j��ͣ�& k_��8�RX�@�(�G�7�1�LY) �oͅ�Ԭ��ʭp�R��Ҹe�=��G�nu��k��8��Z�bv��
J����-��MyS �����υ�� �z�X�܋��p�@������u{�6�h/�<�b��:��V+6dL�s���W��x)�Q�L�r�3��:Sڵ���U�������e`�4�������,��,�_�?�b� Q8��3�,��"����� ���jF0;E�q!O���aѧ�n�"l�O�R��%Ӑ	�|�Z�T����o��_�-τ�>yGi8�v����[	�|�YPa�k0"�Y#o��C�*��s�hg$��2�KE|a�I��]kCR dЄ�X�� ����C�%r��_��F�y�N������ߙq�y<ѧ!����TC�K��{0l�ɜ�}�}1ސD�}���.����́�MK?r:}:�vph��{�$���	%O"�'���{�PXڭK��_���H�Ԁ�0	�thtҏ��f�	�;�xq4�\��e_��'.�z�j9t}���X2j�Z8����j��&��ew�?fP�W���&�n��� ^�O���BT�G��M"z;��$ ���X�*)��pi���eQ���d
4u��}��q�H�c��F����3S:%�إ��M�^��V̮mӤ���N���Wh
�[�D5­[��!��?ΖS�d�nK�'�Ty����&<�3ꍢFꝶ|�8-;Q:�M��������A73�����6���	[�X�o���fy��%������u Y���
k���)QtN����7�O|�3����i��BT�<P^���'�e�-�{��E�#w�Ȧ˗V��>����r�}4�q,�	E�J6��*���T�E��i���a[�1z�8��^��H!}O�pn���(�v��
px}�,���y]�+��c�E\��Uǡ��C��a�4�ꘄ#� ra\ݨ��"�H���4���L�R�]�i��}*�\2nhq6���eh$�+Liv�J��8B���@�D���p9��S�b\��i�uP�+�j2�Y_X� .�����ʌ������s�?XY]��16#Z���-Bo�k^fW!%�m�������p�G��>JWj��+����++j3�[Td=�j���C/��f)lU#j�?���G��¿� �dqj���?� ���I�7��R���>F�k!L��̶�^�{A��`����j�K�m�����jka�	V?55���`������/���|#:��� ��)�8v�W~�!�&43u u�Q�6�:~p�0�fk�j�9^޶c��_�R��l+�<w�`��(}VB�7�8	C�{XH�S�������g����%- ��r���X`wbp+��nf"��$]��0;�g>V��������(��c�F;(֑�b�f�F��/���+[����-��^��kE�h
�@�t� 0语Y;���sZ��>1Ϋ�Y��T�	G�Q�����跤!��Y㉿w^MF`�3�]A�ƚ��)!ܫe��8�B�扒 ��'��j�<��0fg�N�����Ζ���eo�k��	�qO<�	��Ӭ�y��F�`c����)�����=�GX$~I>�O�;���7����ȇk�������C��EJ������U���}B�����R���;��7~�9?�%��~��^�F��A�<p�Kb��i)h��k(}{�m�n������l�������������Q�on��⟵N�
����0$hS�>_&�jm���\|�ь���p���3�i$#4p�,��=g�����.[���[Uy�G� �~Tv��6��p�Wu�#�G�D#MK�Ny�N�M��t��7x�����Wޘ2��Ɗ>�֔@�\�M�N������������a"v(j��!�7h!�$���e��b�|EE����H���3H3�k�-I�ӼDU�����P�L|�