��/  ��E騦�B%:��ي��^���L��G��|�3��F����vB_L���H����X@�&f�a���G�F�j����[����ˉGυ�
�ae�"AE�־Ϊ@�I��s=T�z��q��'S��G2Z����>����'�7���GFި̻ޘ���8�E�U�Hf��l,`x�5���=�?�������ٱ�܇b�Ą�(W�h��\@����|ɴ�H]�j���
�#1�S影���f)���j�Z��}�W��C�H|%L���U�	~˶����x5��Rb��J��p����'���˲ߩhz0N�,eQi�x��r�uc�>rs������W��I���>6���L��S/*{�Ř^a���?����<�J�Iy�ͼ�3�
���3���w�x�׫j�ᇟڙ\�W����;�Ҟ0�fl1/G��� 9`�D��557	��	���G��"w����h���uqd	���*j��#6��X����#�Q��󎙺]�Z�>�o_�
�(�h^V�rЌ����~v �[s�����W5Qx���#��3��#��H���5���*��i��nZ�{�`�����:U.l>g:�b"�C��3cF�r0�|�M���yㇽ�����Rd����N��Į+���79OՐ~�Wl7n� ."�Ѷ_
A)�J �:t��Nǰ!�����\5��$���Y��?*N����F��=E9��:w���в��VZr"g�x^���b����t��ޮW��MЃ��ner>}��}>�H��m�KR�v�JB8��fѼIp���un�S$���Id�����l^�G�Q�0mL�ß?iU����F*�;^�ERg��\~ fܾ�`�"W
0���At+�<�R4 ��J���[>Pσ�Tp�g����Q�,���zɃ;��=�f�M��x��=
��Ph�E����
���5B;�V��Ś����P�(Ӂo��%&�kی�s��w��it��7�O�e��b8Hgm��>���Rk$�n�B�Y��h�����/C�(��SO���v/ꇬG ���]b¦���a��yŨ�M��G������|E��,ƦO��\�lm�"�Zee�ci�t!��2~0��[�NeȾ����܂<�̸_��֕�eV�QTq�������[���hv���T%ͪ(��'�5���������@���xomZ4q�,�ݳ�\��;��|f@�:}��2u���Spn�x����v9�����=��a#+�H�*wu��@���Rvj��(�e�}(7~���Rӷ�^8��R���3p��-���Q%BmH�׫��� �����q�-��e>B��<d�-NU
�����:�8�����ӻ�9�}/Y�D�0Iq|G�����'{	����4�k>��9P�6���v�]��],�黉:�`�4oI�X��lOu�D�܋�;���.,g�Z�[im8�:�t�����o�#{��&�X*(��bH��V�L��G;8��ٲ ſ�i�kf�"�bPv�R�+�z�#.fh�vsKʙa��(*@È���w>I�:��%���&V��ދ�h�4���'��L2�-�`~�� �~�f�yĢR��H]��W��2�cg�Zl��5�=Wsx��*���5�~g��3<y����+v�K���!/m˨�TNf��yc �������.V�����/8��h�t3G<MA��K�W��֌��)�'pGn������X��Qwq�A`'�*W��-������=���c��w�B���2��4e�T	c�٬���~\)��,�9�J�S<�y�L�+�Qb>?1���i�ء@e�z�ȡ�u�*�^Ջ(!�|�4�⊞�F��>s-m��m�K��A*�j��/�M���W�޵	�f���:U~�h��9�M�,��jŝÐ�5,�O|�Ua���2-@Q9�V(F�;�զ�B�J0.$L�쌬C �S�C�;M�n�r�5.'���k���d����R�J�Vh٬v���5�<PE�[��؏ꞿ(�B����"���,���b��R�6"'=���9���L�B�)��u��	��9!��y�Q]�ǎ[&i�|6Z}�=o��,�[�*�s���{:k}d�<LN�����\	��HN�b���6d)0����>ƀ��p��ix���p�r��F�b��p�]�.�k#�]�PD�B��"��wĭ���(g��8��k����<��E�ͤip͏��>x�q�z�46�e�ЫP�W¬]��|��&8i.5ҹ��3(�8��N����i�,��+�ԝ��x�^�?���P���{蘀� �+���
"�c�D�
 xr �L����*r柤o���_AP���\r�����7@:.�����x�1��Ҥ�k��������;�����+p�o˹:��#~�ٚ�4ҩ�f��P��N&8�H`���Hޟ����.��	���`�#�� �v=�3Q�k Yj�'*V7K�,�-��O,��FE~_EG�N���_�|�� ����`4�h\�J��� KҤ�z<̶�&�U4��#�4G�r�k�=�sdA.�.D �E�	���/�D�~�oS/�`J�-�������p�3>n���T�����$o3P�jM>;U�ВM�
��]�E�;#C�g�GX�	O@����:���`*�u����ߊ�r�Q=u���7�@�N�?��v�we�ATS�J��E�`�R%m��<�	k~-��B��ă���#�������u4z)�4x�Z�IJ�t�s����NMP	彭D���/�m�禠�\8F�↑�����,E:)D�1� ߇}�\ua.�&w��E�#�m�D�H�