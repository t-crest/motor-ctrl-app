��/  ���s�*%mŶ+ln�W�L).(	���ĸJ����� ���[��M��|�����BɼP��7=¼I7D�ONy<�_�'1��:nZ�g|��ӵ=��k<;�����TT���<ɱX��|:���{L:��UY9Y{0��rPOSkvL���EF���"�`/V^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK h)h-^�z7��p�q/]%��Bt�e�w�>�/q=R�t7~����E�fjZ>�V;��A��BSTt��4Y��]��+o(���]b[�p�NLr�c��*��͇��w���F��6��>��s!l��'����<Z>X�8���&�D��4���S���FzU�U�$�J�����5ԀD���G�z��o
Cؘ��6.Č�.~j�@f]CaU}��C-5�ɱ��_��б<�g��ge�,�͚@ﯵ��i�g�x%�^f5�ڎ)
�稘f�V_���n�0+=�yn�u[��E4U�k�&��ȽϠ�����M�}u�=M[�n�^��R���#5qb��n�M-� j����1��b�9'�G�{	D�V�t[�Ԯ(x��|�h�6�;&`O�!)��p���rQ�كb�� �A6��Cu����D��@��y��p	b�����>�q��D�e7I�ɧ�W��Tӥ��qhр�ׄ"��4����{��t|�TP�(�7�!��QK��Ga���'�g�z~�l�soUaW�V���x]l)!`'�v��%�V��B'�*ֱt"���ꬑ�Ǧ�W(��Y/~�'�*������윐�E�V�?�#p�d�gb� �z�a@(h���@h/�
��y@^h�A˻|�ps[!*���Sn�
n�$��K��5��)[���[ �G�j��:���W�/f`�?n�b�e�`N$����}@�����#���Ϭ#�Ox�׈�5 �g����2.�s��6P ����Z��5A����G� 1��*T�ȾȰ:�`	t�Z�ӶGy�ӠWo6���۠=��H�e��m$B���Y��y0��9]-�㧃��t�l��ziq7E:���G�H��`���p:��g�ޥ1�ɸ`�W Cc��D���]��Wϖ��r�f�w�O}�te�X��
�L�W'����ޡ�u�Z->Wӎ��--�N�8�^�;0w���k�k����>ߛ6dH������j�E#ئX�8if�{��+��A�D�'��N��)�BBڏK�i��z�f5+�l0
�j�1_x�DO$wwU�ʦX�؛������>�/a��]��X���0r	��f����گ�㐮�����^$<�p�H��o(�#^�Ĝ�H����`�K�00�Z)�˛E��*��ӳH���o��I`d]�Ϭ#m	�)_P������GhP-clV>�W��zI��?��cZ`%8>�;�Ę!����� �3�I>3<��z�6�r:be��
���5=�o�߶��C�D^n���Z��K$��k�p~��;+��0G�nka�a<͝�SsVL�S{�Gʗ��ǈ�Y�5��j���r�lF��*!�Y![Η;OR��g���:1J�ܔ�����᠒sq3v���G�Ʒ�ڛȕ��9Šܴ�8c26?4q~x_&vS�M��@=B�/6T��vM�|�n���Ȁ��߲n�u\���7�.Zݖ�ۄd/�h���2Ȏ3)�"#o��ъYj�WR�QH�myb�F4O�Y�Ȩ �[\������p�lj��Pz��XL��ſ�1��
��p�1��$#�-�%�Ӯ��p5m��ҘTf�S�1h����� i�As^��.@��Y��p�V�w}h>�{�Q��ğz¿�③M|���|f\��mw@���Z;�}�Q	�]��(� �C,��u��h��F7��r�n�q/�>x]�5�ӰD�S�e��m�6�s�L>i3��,�cF�ݍKu�Nu4-��|)x>H�C( �Ђ��BU��O�Lr+�z�ti��&���.T���x �=h��7}H��x�m�̮�2�L��K���ͯ��G��xˤ��QW\6���43��G�����W�+�`���7����>����#�=�6�Zr&F1�KyP<�9����(Z�V��P��9IJE��QVK:���KkgH,!¨Hbj�\��;V�/��څokZo�<���~����v��ȴ1kL
��&@�P�-r��T�ǉVg7��5CG�P�w�Xq����{3�N���u��� ?�S$;|�u" 06��ǈV-U�{� Z�� Y���B��$x�0]ZgG�W}U�7y_��F���W���;$��U�'{.���|3��������.�x�T��
{��ɷE۹��=����@Jw�RyvOp���	tڔ��2[:a�r�0�tves;���P�N��<x9CA^�:�T���,Ƒ�#���ݻo [��E��}��k��d�U���v��x
�j���>�>��ꓪ�A��Rd��c�agO��YXl�9 c"�GA�[w5!C�
J1�,��n��v6qPv��/���&X��,�3�#�@�6<fZ�A�y{y7� ��X.wd�]��<j��h��`�ͥ�!�����s�̼w��ǚ\`�B�Hb��C+,`B�^�����G��AA�����]���c�d�����$;U��`�ߋ���	��B����5�5D�7����L�� AB���ΞPoh�(Q����4��8���C��	p
����^�@95ַX���)�?�I�]��zV�r#�-P���Ś ���4z���9a;��E����jUo[q�S<#0�޺}��G��
{'S�x/��:�d�p��}��g��R��x늝F�}����+砣����h��1�4 c-f��]g�{1�=8v��<�FqD�~�T�X����,𷢈�܂�1�«����%��,�<�	�_���ƺ��$�nwR/�{���Q?�l�V`��v"Á�6ș(Ϊ�KIH�8p>M{͑Vo�_r*%Qf��;�ӄ�'r��(�cV
���d�����u�B� �9���5Yʇ��D�Jo
ǋ��N�j��6g1����]<J���˹�5���~r}x�؊�] �\e���'�JѭiSC��,{  Th�S��Cti����F�ł��8��r�'�q:�1V4�35�c��k�Z����e��e�#ս�����;��5{_HQ�[��-:�;`eH�]�|�=��}��[��N�
w����eX^Ӊק 0΢ ~"1��<!5�)��R���U��Y Uq�mԠP�9�qI烴	��~ޭ����+2PD�����y\�(�ď�mi��y�������p�Y ]���-BV����wE��C=P<&�T]�R��e����^C�Di� �� �֜�J2%o[/�
.����R��ٱ���XX^���]W��*H��tLL4rTC����u0����y½5���2Oӥ��󪕨zɋ�� Uڸ�U(�h�-7k-ɒ!�7�ϵ��ԇB]X�^�c��SE�j�|�r��;��9Z\_�L�o������ސ��}
�).NQ��jlo���� �t�К�/g�z�|вt!�Vgf���9Í�й�7�!����b�	���	��5��JvM��A���GNXmɡp�q�Rbה�Ւ�'��-�?"�nm2B]�n�+��L.�H
ś �_H	��.Y�5�#�|���ZG}J�4��ls��!"�|H_�N�n�Q���t�U�YX��ڱ (�J\[Z"=-��Yf� �4���+D��x*e62�����vF�| ���T�� ʧRK��"uf���l�P/�}v�3�:�)�]՚:��Y2�O����@��K�'�9Z�qI+5h���+�{�vX:���ܔ9��V�*�}DW?�e�3���fu	��D��$��*t�����k�U�!��4.���v�f�N�k7}[�lL�����8�\�]}����׶)�?*w�\7(ƍA����n�Φ�3O^���c�����R���v(�]i�>��t(Y0<�(uͿ�bSm����*(�o� ��Ɠa��o/�=E���1�O��f�)���cZ=C�x��>1�����J2j���fO=�Uj��@��wƹ�P�M�W��*�n��:�X�?Ěj�\ezb�A��v��ňH��	�o��վf��/���?=����=`�೺��L�*�K��S��l�K�
�7�Et�l`�L�s��c��x<�j{pU'�R���Bg�0� �w�5D��O5,��1�X��EZv�H�����X+�mWG���jEw�;E(ryj����yT�1/�� J6�̷f�~*n4�"*@��ydjP��<�2z�D�*���V����#��@��ۛ��|�9�2���qBz͇F.�j��Ȗ��H|�X#e���i}8J�������J���|�n�T�=l�x>S;P�7�eW��bc*���f6z�		K�T?h��n�t�S�V&.�Ҽ�����}ި�X�.":D������$,e�Y��\(K2��Q�_pd3����m��_��t�\�~���(�^��w�w�2s"s�F������m=EIg72��3��:tO���3_Rm�RٌղeXE�4V6�8�\K�a:�T��T�J�cnW����W2��d�ݲ-ge��|�@K�A�tj^͐��-P��L\�����Ɵ�)����ID��Ǟ���v�����,���pEr���e�A�<����W^�0���������ӄ)u0�z����Qij�;���@+���0ׁru^�p��^%L㡦�H�@�KeU���q��#�"VS���I�Y�E`m��ׁ�G4w$q��93��n������$T�:Au�Bh�`��V}|8H���VtAZ{N0"�u�y�T��3�R��i�HB�h�0����R��aP��sV��B��q4���J��w��2�$����̍^q�Ŀ��ؕ�06Fb(ad���<S��Q%�n��m���1��|�6�b��{~�hV���Z�����"��+�ƜA����e�͈Xt]��=�C��X�*�m.̾�8�&8�DG�/�D���0��K�$�a���8��}��͊r��Q҈�F~�)ǡ?�� ��)t��+l�<x�:La���Z�۩g`0ւ� Ϊ۩��.T�h�����i��<��"{JE{�.�D��o�"��	�]�uo"�ג�Ƥ��"b e$��t�y/��-�0���O�m��pҊ�����,�8(��T�T���׊�#�N\B,/'@��Z����S v-7�n�SC�{�|�/"��.��m*qQ�*N��x�3����J��'k�f%����-�b�׳5�(��V�-3��U3`K��.%r���`Ϛ��cU$�� ���Ht-�滸"��-6s+{���Aj�� H�r�M����6�X#'�2+�T�^Pg�U�j$vry� 
���ֱ�v�!�z~eX˖�l`�C����qu3Q�!����H1^ɰ�TKj��մ���D���tsJ�f�Z�d�#�GgN�#�b��ۻ�v?,��~�GZC/w4��An�@�
�J=A��v��?�), {����Hz��#,��x^A�Q����F��QrYi�(�������&�͠�O��iK�/��ln4N�<Uj�BtT�]���O;����6ZKH7z(<��g���mG�l��p\��q}ӡ��'���BI3���b@��	@����F��@��-�om�r��,�!	�
|�ML
������!�f�?�]5����uD��*̯a��i��u���0�	S�!���#nÙ�ȣ�.�I\��`!���+x��A�;ƻEs�u{ز����YI�ߩkCa��Hʶ=�w}B:AX�UA�s�)�9�d�1� ����U���D� ��Lψ�Y�N\E��v�-�~�k��T0tvvjugm�
1C�%bG��n� ��#�K�uA�D��ᕉ�`Q'B�����Ng���R��g_�Pڜ������þ~���u�ky�ԇ1��Ee�]��Y>���҆��{Y7kXI�B,��W�8�2�N_�D�7��q��W��� �f�Ӫq�T�+<�=<�wD�_���6��[b1C�@tM�ϯ|�iE#"�f��������Z(�&�y����c=�o�_?Y���Fb�d34Y�����km�UBkR�4J���P����2�0�5wn�����?���˛��S�~��#�v��UV���*��͍xR�D��_KqH�;ngT��>�~�1�!�"��k͐�#�#G���6§d��Y~�P"�ն��O���P�CiۇA8h%dY�/�RU�?�ǟ����@��5�����"Dz�o�����-qǛ�]���^�뀟�\_���=;�cT6|��9�@K� p� ���Q�o�+�;�у+�!¡�	����!�Ob�EE��Xq�iB��	�j�gn�=꒦�� z!e<��Ȩ5h�`5RW��*�i)]Q ��>k��	b��q5�z����ì����[�B"�֓=Z�r��Rr��ߤ(S⎪_yO�r��Lܬ�h� "���\%�M׋0]�S:���ڮ�p���.��-T�l���۟)��0H~H�+��>^g�������Nw�Z��R���h�S��Ire'�S��=N����mUb�Ǥ�x%�W���J���]��3+L9_kh�3уԼQQM��,�[�<U��cy���Y��}>eYHx{Z�o�r���?�J��dΚ��2�ӗ�v�K%����F���3��"'����?j�*w�v��w����Ҡ� �
�G6������@�I�y02�k(L�]a-�."Ӻ
�0r�$c��p%�,JGN?�_�r���|���LP����P�[���J�%f?��n+�ՠ?M�uI&��0��?ǔX΋yp
�TeV�e�쾥��]*�PJ��~�<����x��z�����yu�E����I�e��y#O�0RQ��0���<�	�%�O��5�,r3f>[T����2r�6K�/���ؐ��;ʴ�S?(b�4Z'��3���#�x5��u���V �A��AN�dwc/�/m��1Pq����p��n~Y�x���=lj��y��9]�-���$��3ĭN�2����u!Ά�6̹��a���E�Z���!��7���,��/�#�1��"��J����.�g�Q������2�E{�?�s3e��1q�� �{G�<<�VtE�m,	Đ�"}�Ӟ��~��\*�ڿUN���璬}�E���ە�4�5o��jnT�]����A�k������s�9�����ko��i��a��8HF��$;���%�r�}��F� �-�(YG��K�Y59���.E�Q4}ƫ�}�����>��[�n�*톑�"U�U`4fg�.��L���.f����7�RG��'�.Dl�eB�^c*S�V�C�mo�<s���tϛk%X�Kr�>aE�!���ƕ7T�t�TQ���^�d^��'����.:�*�vH�"���w6&�"JP�d;w�%n|xy��i�
܅���������M�EQ��U�nh�f !@C�S�5w����{Y�A�i�����:�[n��u�z�!8��.4��$�`n>��M���wH�ZO�XtP�V��G]���j~��$Gr���}����Z\�d�r13~�+[Oຈ3��d�O��'*��K�Q�ܴ�7\���ir���̰���.��x��<����^��<��+�C?^*�q�:.\6C�k>��cV�aw�[
���F�|Ղ���\x?n�s��,��Q��Z-YMv���`�rO2-�3�8E�/���u�۱*V]%�Q���Y%.7Xʓf ��n��L����K�ˡ[���d� ϻ
g��y��+Z������ÜET���/�������?|k
8�v̤  䓔Jc�r�m�l-��'��j�V�������NJ�R(�������J�*ݝz&b�
�U��	��]��R"�ݯe>�+���O:[H!Wo��ַ�Q��,
X�}��r�'6�/�ޙ�uA�*6pK��b�$�m�A5�
Qrk�j�K�2E��/MA�w��}��i�Ƒ�N:]drM��Ɠ����8Zuc	|�4��V�P�� 5��.�X)3k��ꗊ$4>����2(��-��a��HJ�z���~.����ك�a@�ȱ={���㒟N�����*����e���#3k�z+$��bٶ�'֋�J��ˣ�/����Ҵb����ӑܞ�hB��ܥ�����6V���d��זHBnQ����m�E���YFe�+��P��]��d.�nB'�D�H���5��79G}4/=B?vٱC�i=z��~��sP0���� �?�̉zm�E~�P��cB��[T�4G?B���s�2Y����/?�5�1w2�\ ����!P}}{��I��lH۵��(v�3=�#�$G&<֘����%����r)Zu�VT�b���t;��Qi����f��9���ٹ��1�m�AL���LL����sl��|gX��5I�=by�KH�j�#���e����1}��t����^a�5��ǩ#��R��/wL֚�ju�E�Lڟ%�v T�B�E1?�0���s���o��(���G��xL�t�W�����A��d��m,#λT�n��4ϵr��V̲�L	�R{&8Z.��=)�՟�xe�������:d��B���z�֌��a(�}w��i��{0�쬋�s~�:LĠ_)N��S����:�-��cm�.Џ%s���G�>dN����թJ|�W�ξW�>�w2��kiv�k��n �w
5���ƪW&A� �3睷�/xv�v�<��uN$�Կ�u,�?-'��O�U	{���a�Ɉ��\�v:c�W�SI&VƘ�X�a�'K�. ��z�oq�_�U^t�xe��}5t[!S|��V��,r�˔��ҧ ��c|$�#���]2��BE���t<�g�;s-Z�{,D7�*&Я�)WJ��'m*�	y 
bP���O7�J�Em�@���:�.����l�J΢���=�v#S�d�y{Y䲟'R/+�9%�g��P��Q�=q����A�@:gp��-ݱ��b��O���qi��<�/
������x��11%s!��G���ηJG�"�K����DA ��x(��o*l-)`��㨡5Q;$�A(�
�-:y�QȬ����fR �����p<]���(a�7�iP?^Ă��%#	���,�p�6?<_����ǚ������N�瑖�E.z����b
>����q�� ���K?n��%�.e(�9�H���[�gN��D�hC�`Q*��% ���,H!����0�
�^ 5׮H��
���`��}@�D��⪗ ����jٍ�����EE��ݘ|�(U�!�+@u����G󟗗0V[�f:�C7��
�'�� ���d�Z<���YH*#V�Ӥ-6�������n}����=6���K�&Z��۝�JND�4�f�5��q��K����A�d]��B=��BL�F~_�͟u�R,I4h�SKCN�5��Ǝu+2ǅ��	���ğ���<7�J+�x�[���1�F�b�����u��58�?�T}0��9�8�q��4h����C�_��"y�b��{7�����gVc�L�k4�ޒo�Um#Q���f�/7�z|�j����Ӝ�È���+�}x7ّ��i��n-��r���q��1���㸷��a[x�'��i���[ e��fH5�Å�<E���[�Χj.�=��s�>�d:�4��t�:�ԏ�n@`)��j����s�z����7�ް�;a���S�(ur����b�F�,W1�%�~�P�A3�6p�m�;Q!��d���4����ͮ���n�h��.	,,>1�c�y#� }����
'���5عC(�3���шW�+��&}�;�s2
Z���5��(����5�©]�]-�1\@Whz[�ru>�С��M+���v���=�_р����l� �tR�<��o��U�X�2�k�����_��Qr��ݤ�8������]����h�fd޵xv��x�nV/���}S4���T�Ʊ88�U��1A�s*]��H�����-PjP宎̡ҷi<L�x��×��SHL���h111�����|�_����܁�u��ZU���VX#OYQ�t���O�8C����� �����gG��f��Q9��~�������GB��a�>d��53��H���u�>
#��$�V1��&f Yn�H��ȷD�E��^S����̒�:��҅r7��;���
A�0��vg����j�.�;�=���zղ/�\M�ˢ5�7�Ԁ��T,,�llDR��|�3;.	Fք�,�O�oq�O�#���}�o�#�֛D>�JC�<��/x_͛%g�n�O;�^�Q���7�H����_��Ɩ�*��������\n��Ҭ��\�ˉ"k�nLԜՍä<��x�"-��˒����QQ?��/�.�cW=sRz�����5U������0[gqTl ����僲38��C���~��U��w wu�m5Z�b��� |�����
�Tm�`5�D���Z�w�l���-��ʛ��^��V�0I�ë���]�R�d�$�]�c�h��V�> �md��h�^R�0ck�~
�����j��ۮ(��`�s"@�
�g  ���)4g[�\���ŋ��=��X���4�Ug�C��]JK�7�$;�*�-(Ԉp����0����s�y|d�|z��3�v��q�����˙�kF�"I�`G�.�*�_��E-�Js&�4V"���d1��t�%_a����$$��e������rf
g����a"L�"C
&�B�$�¼-��+�� Z��5���y,�Jim�T�f3�Ne6��?b���HWQ��d�}R�r9�E�ȯ��%�	*@�͛�	���;��gd^�
'���6�sn^SV����}�J���@бx'��a~�'s��N�9��!�4�\"�oV���&�5
Q�o.�nR�}|��O �~/�4Lۿd�9t+TC7�l��
�K�"��j�l���j��X��׋�L�Ӆf���Sy���a�yp���>�E��ɑV�7�Ӣ\��x�K�6� �H��
�&����r��1鞲ch$���읳=��$�3v�Q�Ok�6|)����$����"��q8����%�w�3�ݻ4�n��;OUPK�U/
�ǌ����c:�iY�Ct���^xm����i]����R����?Є<٩�d�]$Ջ�Q�x0����Q�0j����u�:�� �E����K��ғ1�}�a�� �/c��{{��a��9'����Y����c��F�'X����T/1n�<�p����ߔ˷ruũWvw���9�pW�/��c�`]e@���^�-j�6A�Y>�Ṙ�vf������ �N��������h4�qd-(oU���b:�A��f�� s���$�Y��1��Y��+fJ���C��Ƹys��o��rk����a���z��:~o$!�A�&��\U�B����W��\��}<#�ǧٜf���$@���HfoZQ�pX��<PQ��c*Ó>���Lgͱ3������ `R�(7��a��^M<�鰃ત�F8_�8w�r/��9;G���$Ae��Zv��vy��u��%c:��%	z��#�ZY��R��)rs�W��L9/�-��1��`Sf]A:h��ͽO�!��T���*�7%Wx����s"^����V!Z��]��aN�5%�}�~<g�Ŵ��~�YRs������Y*o>9�c�vB�d�nx�!k
~�ݴg,R�J�v�X�y��x>ʋm��О��k\���0�u)�I���ADj�@��^�%Tq�J�*|���,w�b<��<PT�a�\�M�0�h�OBy��;���*KJ!"B>:���P��S<p���y�C�`M��El�(�C���|`*M��]��Gx��X�_�q�*9b-K�%Rgl�o�a;B�|����� M�	�L8�I�:�q��q����.�0���!2�7�4�6�cX����CGD���L��~��Ȣ}?��kp�ɘH�ʍV��Ju�W�Q�m��*F(8��ġ��39޳�J첆#}r����� 6����9����w�0�F)H�`��൸��-�b�ǉ�6{�͜�A��q��
w���Z6������t�l��n��9R)�LR�94-�@�i�9���'��-&?<�8x��gvq��ǧ��Ra�B�@��&wtEǨ�j�ó~[�*|.�{�^�f�� ��O�ns����DT���G��7v� *�(��f��1�rgVw�fC��"Yst^7���-�Bt��텉.�C5!d�`���^�(}��(�:���S`���&Z���t���xF�&�j)ת���X����x����Q�f�$�7�g*R"���K$�T/A��2�*"&���ţ�h��(ӵ0���yI��]�'���M@rC� ��EL�æ��o-e���G�i��=-�ͱ��4J�A���RG	b�&*����I;��U�p�$	������~�5��]�L�d�Q����:��oX��/B�������p,Y5�b��O�*)�}[�xW��1�13 ��%���8K%EF�w������}��މH<�X���Җ5к�k,I�i|fgU��ZM߰����6�ǜkR��k˺�