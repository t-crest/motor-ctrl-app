��/  �Ɵ�b��b�o��y<:s�S�I�;��y�F,�#b)���2s�F���$��������	m|8���atl �aJ��]�N��ͽ!˜Zo�|���ꅌ�5G,Tv���`����E��5@�Qo�u�AK����G��T��򔲇�H�����X"7[m�.w�rApX��E��l/�o�3NȽ��oʋ&��B���Oq��Bz��KG8r���F6p[��J����(��2��~�������,�Qp�'۲  4����-�Z��H���g��R�+7^%��Tj�\ý����o!b��:h��0�k��(wϓÇ&1������w�������GW�ޏ��4G�=h�1t�R^���]!����Cg���u;u�
����i̇<w��u0��Z9J�!0E,��{rs�8'��N��̀Z�$�+�;o�إ[�8{)Q{~�`�ޱN��ǂ����uô�͂*^�~x)�KYt�.o�m���)(�mZ�`�D���T���jo�����Ux_�fio8geV:)��+3�(�����;M��"����N�A�!���ہ��i�]�C�a�4��=u�S��T�]�'�1�I�$I�c�6���d���0�O�Co�ƳK�\Kv憉��8c�9*	'nfP���N����Q���vez/D��f����qd����'e+�Eq�\HAAq}�WM��Ӎ�bq�G�����5�6��D!��F)�EŘ�P�����;�I83j}}��X�=�P�ߴV��J/D�v�U�(o�1 �+uw�!�jaP��%Vq�y�pt�z�4)�V@����z��Q8�QD�U���G
)*���e��oGp珃TZ�}y����49��~���sQ����t��C/�M*�C-���B"X޴�G�׹e�j��@�E�A�j-[[h-�� C�˼+�s��
D�z�2vs[!� o�W|Մ����J�γ���n��^�zv1�����Ddo�a�3NL�G�:�j��Rn�+��Z f�������R�,�r�j�jtkS�(�ͧ�����%s�>�d�p�l�����d[aE�1���Xވ��d-�	�6�` m�@uQ#V�0귓r��Bĝ��9�]>�ļ����Bc�q�����7��u[��������W�
x��As��a��q+^�����=C;e>��i�b�B��\��W<���;���k�!����O�z�q#b��7�NM��ޮ���:Z�F�n�?������_[۠=$b���̓����_���'�e�����X�_�KaO���j��Ɩ4R��ŹqkJ�&�r F��t�G,C�p��O�M���s)�R��qtى��Z������ ��z�����>%��j�И&��^7��n���&�Qp�L�򶪟��k�%�O��ܬrX<yUL�[\�J=�@�6D����W�J7�``�Lgc:1u�fֱ�10Vw�ڍ���G���ص�W}k��Y��zW?�/����Z*G^�e!��cM�3cnt�9���L���2&�'��af�0�&���Ѣp�12 �~L���闤�"V��qX@g?_I�Z���\a�JN*�J�����-�^�#[b�I���K��tKNnK���dGpۖF*d��k�1!�nd	#ʤ�,�-�#P2i���QD�<�.�F��b�[x�^�ПE�QG�����~o��:'�s
a#$uyDZ����Sx��PQ�1u�}��N2�1�84����O{���+ 
�(7��$��o���f�HA�G�0m�̢�C���W Q��"�8�V��N��w����G�PP$�B�l _JA�Q{+����i�"�y�Z���(��gLy��Q�I��Ѽ��\֔
�����
��CQ����Rͬ<��(����]�6Fx@� ��ti8��V��&�����~�A<�mγ8����q���#�R�5��L�Ġ�d�f�4GI�tz�\@Hcm�8UD��˜�ʎ~�/�'0�#�[DS��s'[]��(~�5�o#����[)7&�]5����;Ҷ�~\|��ʹ�~���o���#�Eu��a���j�.�Uv�f�F�W���R6��w�������R!�f0�R���`2�^� j��eo�ܕ�c�em�ܖ�o��e�ܲP��{�$nרUs1��Q��'��N-����A����H�I�v���Cd�H>K��.c���4�D+l:���^�����]��R����t�4!�'��� Π7����AX�PC&��
M�>�Rzu�|�a��iwJ�JU�e�����.9 �(J#4��W�����N��u]/н:��Z�a�
*r���W`i��͚n�WV�(���f��zQ�eW���9��Z�o5����8$'��o��Y�˜ b��{�A�2��=Ӳ;���x��	M����s�c���n�X���[A����K�o��j�>#��1_f�),��;l��� ĩ�ٔ��e7��%�u1Jg��޺�e7���L�Q&@��;��ޞ�,��$`z�h/×�\�\Xv���W��e{�r0�@�J(�L%���U$}�"�O�E����q�����.�.�gX<���;vt��$�Ȕw��s��ƿ ����@�b�2���H!����X��J����־�8����RY��I��:�x*3�ܞ���ǔ�n�*�������,W�[z)�y�FM��G�������ĥ�(=űz���/��E�������d�8�g�F�I�Ty!r8�&Q���g�5uE�Ȇ2ڽ�f�Լ�Jӥ��)֤��ȽP�����5��Z|����Z���>���O��6]߮�O������C5��w�=���Q�F�~��|���`v�-t�fF�/P�N֐>g&����P)�]��� GQE~�W�u^�7�L���!�5I�@�מ�Y�T����J��A	��u�_u��J(�oG1-�|�>�ag$g.Y��yhV9�@�eg�Iۼ"x<��F���O���ȴqk��z#�׏��h�����R�:!�}r��,O_�Tc�+P)��2�}g\;o& ��eO�-�xnV��h�#!uA��7A@�����At[���z�8�����3	�*N4�,�3�a��|R5�F�����eo�<L[xy>-`-�d�t	І�^ܶoPF�����A��H&�m�؄B�ϱI�}	o��һ�������S��r����O@8�����Sq:l���²E��4F%(�XN��>�����(Y!�S#�� �]hb~|e (O˵lR��G��
�	�𞲗��ڏR����`u$��\"�U8�\���XKFa&�c5v�xΈQ񉛓�������?xv�<S���tO\/o�2N:Si����)^Oc�2���,̘��5ӌU�Z��S��Czu
�m��O�y���G��=��$G�d%��4
�,3Q�����3�[#��	�MG��'��R�5�,q��ܟ(=������s[�Ѭ�E~�^�x'�����D	S�zX�LT�sw%�-�T��g�7�����=�m�yGtW�D�Ž$�SCt��s�ɪ�����"�s*�U(�b����VZb��c�z_~�n������F��pt�=�Є��f��)�_��Vig%