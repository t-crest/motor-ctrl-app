��/  ���TCqjN�4���f���X��%x6޸�:^�<D���7䭋�j��]��v��w��äz��|� ���y�Iz��Me	\���42�[�,������j���>����~VW�
�~��DgN������Q\@b���C��Q-�ę�AΓ&g��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<�Rxa?g�j�$���;�=p8���7��r|U�����s���u� (��A䖘n��D�3>�XA9Z��+�w�|��3.w���,�����j]l�j:~Sk�$��E>s^����"�k�-E��k� ���|���XQ�IDr�Ʋ�[��1���]���݇�w$h?��L8¯�����Y=i!e�R$�K.�{n�9ߧ�.�xP:���6��0���_��ȃ�%���Y�V|�g���e~E�W9h�Dǯ�_��,KK��
Ѥ�RlaB�x�Vѫ�w�����A�b�G�)��RFN,/$W�@�<���pM�+g)���d��T��[�i�p���]��V�6��~QN����K	��q>>�o���>R��P=����%^Nz�o���������=ڴ�<�e�/�	������f�8��c{q�1�O�^�U���k�1A�S&�� �(��Ԉ�!�B�2l���+�����g�!Nl+�ʻ�2�������kY����q�;����i�@c�L���	�YCb$]J.���$�["Ч˺<���R��O�@-��Q9+�����ک��vBV5R}(Nd.C.7�z���=��١�Χ�<����9���C�oʚAP���ӂ�	���w]�]�]�J?Gq��ߩ��@�U��*цv�j��[7�S�_���I�8�^��;�p���Iz<�B��$a��i����kQ���b���_o�ݡc& � M�iܕ���ᮚ!�b�eÿ;�Ú)�n�?�nL���X�ȫ2� ��U�Ma�"ț_��
��7�-�z�3G��I^mNG8N�@qq��hj��c�tZj�ӽ�DJHc	���j��Ef�d��Z����=!1M�w�UK0���:.�޴�K��z�}GF@�
��	�Γu� ��G"�^CcgS���k#��6d��i���N�=�LR�x2�\W�]hFO^˩�&�>�/@��m�������zTLf����O$~Ҝ�(�7�_�l��S[Z�l���h�x�&�Kڷ��L/T�BJ%'��0Q@��������XRa�`A~�X�OJŋ�22�[���tR����R�Ǘ#��Y�;��uH���Qj�s�%0��x���Jr��0 ���8+�Q��q���A��J�-��=�U���G3?���J�÷�s��^{h��!w���ǅ� ���A3�ݕ�6��JH�9�n2�u��֢5�y��ϧ�3tY��dn�*��N��z�P��־(w�@f�oNZ�m���4�6}����*.6�°TBb>O�%��dW�h`O�?2KҪ��ؾ��đѬq\s�K!� ޅ��-y�5&XXՠh�٦9���L8��������I�S�thsx4y��db�6l�ў�
�U��h��&�2[��1(}�d20��J��U�~ro�?�R�W�y�gl��fB-� q�P'�����03I��K�v�_���h�
F��J�1�94�������oa�N	}h�g�L��Q�7 m�3_�T��^=�t��S��z�s��B�WJ�X?�ƕϴw���S����N�fڛ�6�֬4v<x�^��q/�(Qg�{L;��؅��y��v�Ro�� t����NOæ}���ge���
^		��6l1�~#\r%#=��z�SD����^�6*��{������K�TD��ۋ5n'�����RC���tt�M�u���o35���iY;�cs_�3�2`�4a9l�����)�a�&��F�4iw�(��5D�"�{G��'�&�^�+!��T�/Bx���3~����R��\�"���A4��������j�ը�4�n��W)u�ㇻ�kIgj�`T{�<\�,����d?
j��P�fR��P7�+,�`�ՊS���7�%���{`l)����;>:E�����˿p�C �Y�&��M�a���=�l��|h��BC(xi�)�l[�x%B�Tm��H=N�� �v*���Ӿ��VR3��"fp�`m0���#�ح��I�����*�v�F5���ʙ����g� ʧGQ<4r�b�v�͓��c��.�^�ؕ(B�����Y��+�u���`"�q����2tf��"Y[uP?�Hn  ��8��H�#�3i��:]��^�z���}��\��D8P��N�5>k�C3WLmO�u�Ѵ)�����u���w���Z���`T��cz�n�-	70#12�W ��S�=�����ut�%��&]d�$Өe����w��<ǧL�M�=ʗW{V/���]����x�6�2e�DY���&3�i%#��3r�+���In�"�?Yf����'��)��Ag �¤��eUo�3��]li��#~͋W�J+�{�	���%k����ҧ�y>-�5�Qʷ�B�Eu�����̀���=i�!�2,� e&��^��kK�3�F�M"�ܙۋj���O�V�p�g:�A��� �GN@��
�H�4�`�cE�B;.��i��8R�lo��ЃԐ/��Y��Qh��zny-I�o
�zsM` �D���$��xS1r1G���"���A�G�F�}��P]��6d(�>���g-�bOD}�Лɼ玂�H�ª��?��Zߩ�p�VH-����.�w��M�eK�"��������JTw
�,�E��֟�X�