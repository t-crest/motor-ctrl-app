��/   z�d|�v��K�6��w�C1o�ό�rq:���װ�`H�۩�5p��p*X�h��ҏ�����G>f&�}4����}Ǎ��S%��TXyf)�drZ�p�%��)��$>*�#��hN���cS�Ւ(@���D!�x�%�妊�2+o&��.��|�^��<�J���6�����֕�]#{��;̔�Rڢj3q�HKTWuޭ���VI��l�ڋz���D��>�,~���j���������>���@`b���W�ɫ �r�9�������R��?c���8����b�lX蠷��d�J�����[R"���V��lbWm�j�r�wKl_�e���q��G�U`�lx;
����?��"�
b�v>FF>�+}�N`�X䔃�c�*�~�mJRt�M�od����V8nQ��i��������\� _=���J�������ǐ��B�����Mn�G�/��*J��Z�����F�y��4�s�S���Kn	W�Nq�zAZu�;z���	u�{G�o���"�4q]��!&=�6��ۤ/Y��M'?�^+����%>Kՙ�7?��b}=���iH&�}��e�f��W^N)Л�.�(�c8;�7���e���n''$���ZV�<H��@Fɥ)Ew0k���m���8��
�l�ŭT�12���@$Y�oO�k!������ ����K�_�?-M>�Z �����d����]o{gU`�w���ڑ.j�A~[�ʛ�r�:��B��(C�j�V���75-W�^��VK��4��SDVP_��[�(�]h�N#$[�Yo`=DI���t1i[N�5!�ͷ����g���ݴ�	�˒�4�T�Ϟ��z�R�L2��m�Qɢ=u�I	�C�h����6��B ��� w��-�,|EV��`�Xw!���P��mվD��qjѤ���e�Kg�%��2fOw��'�<.e��f�.$Z��c��*2ɸ;���E<HX-�V�-����lmk�a!�E�BhP#�����~� ���;x��G��RR�@��9u��m5ײ��LXl�;�@�uJ�Z)Z��m	l&��fj�,�;s&��{)J�9� w���(AJ�wo����Xo���ߥ�`^�ܞr� ��'_����O������-d��K�<��;������$��^W�h��Eq�`A�)���m��I|b� k�n V��h��a��#!��d}���b3��0�q�)�z�9�k���g��{}�a�5d�L?���e��/��w6<�y 
L\��8�l�V)�;�����9˼��BVZ�nt��o�xZF-�g�/XAE�����s2�|���7���lF�9А��<k𡧈 &����J��:~�����_{�,}C�Wn\k��pO�U�C���D�8����y�C�k��n���ƥS�_�����g� �F7��Sq�oO��3q*O@�S��yo��J|�@� cޖ�.n>�&�|�A�e7�؈R�>�RD��R��h_�e� ��̴P4k�I�1��l����|T��09���8Y������=$ �Z��N�R�����H��⾴�P���:����%S��W[Q������k;��Rr�l�L�.__w���M����nH���E�������5�c[�D��C"i=[F9A�d����쯊�12wRY�*�-!�2�AC٪]{���2�j�x�������0�d�z(W���>���Z�r���i�#�o��趿0v(�#��-�p��^*kF��/�������}'V��8�����%�6��*ޛ�s�<;B�is"��ŭ�)���3B��y��SU-;b��I��
1��q�	���@YG�n��Z��&��UD�c����]�L~�&�g���yN�r�:X�̎ݺ�᨜@��X�
dM�r=:��i�s������z������2�n��9ו"�g^J���/�Y�`�8ai�Yn��[�E�R[.�(�����E�l�*�9�پ��<�i]����枱c�ӷw@�������T�
���3�6b�&�z,�ڃ�~�܈U:�ZY�9�q�F<�i��3��|���.D2�M�f��6痚���T��S���"w�����O������D�l�
��$���K{dF��wD�Ff����u�	������0=��.r�?�0������RL��M���y��r��4��Zr,�u�O�h�,)�#�������@iV��
.4A�.��4�r��cIR��!3��Vv��0k*����oƑY���@��<UBY\�TK���d���9��nJ�rN����cM�t�uf���\� &թ�lx����b�\�z�l�`㑥�x%�ݥl�x�<���n�cJ�� �peK,Y����N��7@�y�A#5}���$���-+����`^����OX�4��D�^w��VZ��_^i�����!�3�~�����%�ae�2<���I]���_�c��ZeY �� +��ca+f'
H���D����{��C.G�6
Sx5�Y.§q�X&ʨ9ȼ9m��c6��!�԰l��B�M2���p���_���L^@��qp�>YCO�<�����V��9��Ϻ��b��*��F������&��:c�M�d'��:��"F#>�j%A��%;zdv�Jg��rL���7yiN�;��BH+fz�2�ؗ��e�i6��l<�� ��M�->b�߉n9����^����H3L��{�Ͻ?!%�����v�I�l_����H�/)����(�2���m��n;�����T.+�L���H���������WF�
~pr�[�g�;pN4�*8l {�5Xw<�����L�^	s��~}k��=��٘"�tg��K�{Ho�ț,}��dW���1[�vh�ѠP���O�E�ʼA�rg�w���!�[_M�y2��ν6�Y�ώe<p���Rzs����ow���14���`��M�D�|#�\�5����O7����ae��2������� ��zhxQpc"!�D	��h��-dÚ�ƻ��Ȼgz[���)JS����Ϻj��M�J{��<G^:������1Y��F��z��K���A���FۻRQ���IGw������)r41�;��6&"����kg̸.ѷ�����ag�����j���l�Z_��י,�����\Ig��}�5����2qg�1��z��J��{:G�A'�^��9)��|_87�Ʉ���RS~iR-���\�������'��ʱ6m��UO#}jF~V���ߖ7X�6���w[A�HN�-�j;��7կ��i)>�Z�x)%3���Zі��s2�%���JQ��沏D�ڹ�F�\�H�1�&�l��D�.�$?�W�Ms03�Sr��'�{�ʠ�F�/4f6�7��l7��-�ڻ��<0_��E��'��kH��]	�N��X^~�&ai1����h��ܑ�JUV�������89؀�i�K��a�:����b��,����
��H����� 싈MV�v[I��^g>�=�ŕKg&�e�.gG����R��>����#��N&O���R*���璿�8�d�u��{�yu�;�y�֣������e�ܑ�U�T�ٔp�j�Шė�Y���2��@�PT�=���a"@�v��r���C�T�6ȰB���kkBW���/��L�E�D��hښ������$l���]*@4P��M�x/ɉ����!2��J�)�
��D[��}��YP�j����c:GD�d�2��PS��f�=b!**�sPX�����wwK�'F��3���}qЏ*�[]ۣ��̮V�����	���˧�H�Y�{ﾻմ��Z�"��w0����Z"N��Qȑ\ق/b�
s�»	������H��c�͝�����w)���`W̐�����<���Yq��\̂�k��m�������_�m���T�"j��""��#�֜�ԆG;Xbd�-hTDۭ�/:@5��=3�[�����p�%T#��G���Q�<w~�Q6f0i�#ؼpm�P_"~�s�k�^� 葄�o��$|��!��8ȡ,j�A���+K���;�&�vu�w�PT���aJ��'��v�
c5#���J���Ӗ���4�ni_��S����KG�3��M
ow4vR�B����=2���1Y�f_Y���1�8'�n-U5�Ue��u
�#h5	SR���}`�yW�����4߁�!�a�e� �.)��_0�)-���Zu+��������Z9T�h_�(�!�9G�FɣR�}=��Egg�L~a�R�����"���f���Ҹ%�'8E���@���Ð��A��I��r|	�0�l�?m#E���ұ��<�r�M1Por�D�-��ڼ�m;��{ӥ����@��ē�m����kbZ�����2���+��� ��(�I�P�ҩ��4��嫵mW�Ȋ`�l��?�F0�C���_�0��U܇$(3lM[l�h�}=B��`[5���N�9���6'��q[��n��:f��Sy7�(��C8r��eQm���Ӆ`ʴ�1/�Q[���c�>P�h��D���ɤ���k� q�{
/ib`hA�+�D3��q�H�����{�e0ȅ�����+�vg�Q��4W�X�[Rv�-�UG1!�&�Ls��_�����r�mlslP����b��N�v���2
ke{܀���q���]��D����e^2F�rY��t�Scq��-F���C��ޜ���K��� 6J�W�-�Mb��o��IF"���qQu� Mp��t�~]�/*��x���w��vgg%j�Q�;�G<G�gcM�K=03b��*NY��K#"�:�W���I�z�[�R�/�ژ�no�,��QO���3��z��+�;Fi���O�K���|kt˛#P�*4���o���f���ɦw��ũ�m�Q��L�"�ܞ'D�U�:G��m�}pa웆��SUi�{��#�O���D��}#���ml�xv&$֡�h�b�3�=�3�Ob�'�(�k�sy%̝��f ����9�����*�����^�딭��n[�$҉���EH��W��gc?���qĝ�&����p�L,,370�"��&����q��_t$�������L���ʀ/$�}��a�O'�層�%˜0�4T�%H�\�V�7�\�IC���2�&}�8�KR���#�^�c�aq&�����M�Ɛ7>!^:��0ڒ݆����5Tly#�)��T�}����F��1
�J)��v�ތ�9#54e�},���>��/P�0�K�a~�mX������PhW��J�q����u���$k�Qlg�D�ɞ]�+�f5���)��y��z�&�_��6�Ģ�1����s.� ���D���@�I�๿xO�_��NFP-�K]�Vk"�V�z�2t"��o$��a�q��`*T_.J���6�pT`hπ���l��)1ZC �J}��$K��;��E
��ϮW�y����-G�KH�_��֕0�0*ҍIrdQ��a����N�|g��|87*�M���d�a�v�>z1����6��߇Ck�<�2j�Ȃ\p	jvF����kX����Y� �9l��9/�|՜+��ޙ12<�2η��	���������Z�pU>�Pe=ڡz4)��q�7�Su���'��X�x�r�?V^5\[*�f�?���;��������� �?�1J�U,�Y�#@hi{��-1"?B�[ZgQ�������I1�qU���/��z��w=��z�e��`{Y�I1G����R�J��VT�i�4_q�x��� h7˥�XDR\��T!�����T�yE�h�3�k>mnz����C�t�n.uc�}1k��A�YS���Uc�m/8b�Ġ�s�M2-Q��N�)��[��0�u�z,�z�f��Im�"Xnn��f��4�O��α��f�&
Gf��z8��Y���^D�x��q�q�-���3��q�����=U>�\�:�u�����T��v�M#�W��_bG�SX�!	H�Z��~^�S8���JcG#;�o�!�#� #��,�B�g:��K�A56q ]��/ƛs�ȏ}��(Lt�IQ�^<~#�@��}�4��ey���͊ rfCOe	��K$�0��"
0(Z5FK>��񡏡��C@����ƚ�'i¾m;��#ɖ_�p�@J��_� �n���vh�\�#�1�w)b"=�XGTZM��[L.�}M�z�~�$ix����5v��D�p�-|���g�(-�<���ٷV��,��y�o���'jBE��@⨇�e��$�i�$���%z��i��.轅=��k���֮���9sx׼i��JR��Lv2���(��g���+�
U��s�tJ��jc�&贻+�NI�'���U�N*6��i0�S�/�H"�t:��3� D��Z ��c�GJ-��̶��P�L�0�qF)��zj��c�ބ��8Ӆ�q��Fg�dsC9��bvR��'�b����ݹ�����2�k���ڵ�D�/�ɫ1 �(\�n�XhZU�,�­�mυ�>oH���dP�5Р��	�?(�-'�ǚN���k�;�-tqbG�!.��Ͽ����
�a/�˃=* ��4p��Cg�+���X$���������E�i�|���d�wJ��SN�ǋ�Um��@-��6=e�3�#���^lH6���!��-��'<�3��I��SJ��z�����N�wܢ��(��P���ϾT�<����.\��ߺu���cx:��w�l
�}�up����9-�J_�G*G��@� �G4�d#�ʶI%B��v���~q�pGG1�/L:a:��r�ڮ���E#��'�}��qKw��`F�0�|ECE��[��s���1�.�����2�>�ʆ�A �ڊb�����!����ȅxTe�%K�^��5� \9+A��H�cP���
��kM�upu�h8��4�K������nVc�&�E�řj��c)�v#*�`��<<�=0Cс��W?4�.M�TP���_��<��'V���l�VU�໌̀'��%��t9��M鼻�1�Fb��b��s�ݻm(�
�$&�; aa1>�v�Z���_��T�'L�,u�t��l�.�l���h�Ȇ�Ο\Z$Q�P�w���RQ�R��p%m7:��O�)�[�W�3%YM݌��5�k������1�Y�~����w��z�W@N����ߴ�f��⛹�J��&^��HZ�����oJ}-���/|Ϭ>���H)�!���|�)�ꂹ���|W�k)���T�Ҹ����b�*Y�]���Pk6>� �1��|]�J��F�5�O��8���~,��эg�u�����x�)tQ���u,OӃ�7�&�]Z�XPn�üN���e_�:[Q��P��n,���a�2j�z�H��S%l[�\�l$t:�͆�F�q5,ؽ��F��=���ʅ�f.ݤ���F�!�YO�r������k�3�g%� 7�ʳ��%�R�8mr�T^���_(��@(N�a$�=������A��'��:$}����޴][t6d"����9������,Fx��8u��_��=���[AJ
�6j�]�	�^�����9#�X��c�2�[%��<��#%��;r����a�13�}��M���6�H����Q��T�bҢ�#:3W�	n�}@L��Y��C�Z�y�Vf
�{�PvM.�L<�nJ��I&z�x���͓��_w|�{���1�7ϡʧ�|���%co8|ha�B��`K��|��%�C����Ծ��o�'&\ݐѲ���%Q-��<�)�����0�w�m$:�HQM�k��:��,������$�s�[��Ao��%I��=��`(�@�d��J��]k]�y,�q�2U�T�?�}����χ�I���?s?����ӣ8��N.��u"�~ilݙ�\�˳��z�ī��-�l�D��=�Ƿ_hY<�R�lY�#D>y�|��˔��#&^���v�|{=������Y0���
t���}�Im�TldP�I�W5]��P�ղ�r�n�W��`H��xHW0H\�2�j��9c
����������3��}/�_p3 �Q<rB����5@���@��"�b��b�'0o&��/���O`P�C���E��O鳜�V�q�V�|�r��3�N	�dѾu@aTԉ<���E0 Z��yy�=�����q���t���K�|"�W4z2_@��j����W+�H�z�΢;����w=���?���췳0Ȟ�g��˅k�<xm(��-�4�17���@T���? n��`� �|��Ŵ鯖�E��=aB�~���E�y�~\��^� ~?��a0��J�����ə���ܭ���*�L�a�{xa�x�"b�k�p�.t@9�|-Z������~G�$�Gh/�N�:~�N�`�~�@���� ={ؐq!��G	 �y�@h��v��5g�����N J��8��EQ��ֳ'jWſ�N�����'_�
��yĬ(\�c�
y��݌�J C꛲^�l26�`��>�&�.E�=��˷�{L��m��f�6P��<�3(��
Õ���:ˎ8�3BOJ��ɐ��]y�ʆbRARy"�ER۸�	�G?q����©g}��y�.ڢ3�
�h�U�Eq�[d�B�;k0�0+�Y-����0�j-��"_�,�@A#0]΃��EK+IV�e���QGG����6S�jQ �*��@��\1�G�#Xφ�9����E:DW���k;�7Nc�E���z�4R��n�z]��ZX��u
q��(��lUئw�j���&��9VN[������Bxf���/��]��"�t�YQ��l�]�����1��7%��>�՟���%+���[�髟���ǷᜧO��<�H�
T���ȝFz��돁��t�,�7��|	��l�'���Y��w�#�\&5�V�᫑jl�����R:?֓�6��<ԓ:�&l����S<��A���G�Qꐑ2���_�[��B����zSXBE�����(	q��HA}Zc����� ���*po8
�ڍɗ�WШ�-���"UK\���ʸ�^�O�C�28�c����p�n��q��s��L���Q�������\���Q��~E�u�N��^�nA�����g��X+"%�E{�Ϸ2���(g�~.�"�<��Zn�}���z��ʝ�a����|j�iL"-I�r���SE^b�?���,L�t7Ṗ��ɂY��� ����t�EJ�2���[�.�'��w�4����c�Y��;��܎���K�n*�k�����а�SI/P��#V��}�2���O	�}I��4oe��L�W��^2"��g�d[�M�`ϴ�a�s����"���X��g,�P�*�W�Dy�Zw���Qr��~j=-�' >��̭[en�&�a0�����$�?�/�-��ٿ�6,��ή�t���i��#��9��7�8���y���=؋�DYgAɽ��o��zc�|��dƀ	wהh�a���u';`�ݿp�ڈ�=�VE��Wn��g����aZ^��V�c]��.�a:W(���@$w�:!p�b�d$JZ����ڷk"�˧����lW'��@���5�{e�!��D�)�Y�]�%x�u0�*�Wu�O1����OTH&^����Ht�"�:3<O!Á��=����*�_� ?�Փ�q$��<T���cZ�D�� �yxщ��V������oV���-��}�����I6��� ��=��$�X?�
\�?�LC�͜��w����IF�-H,|��������B��X�
��q�ƕ�Y�R�B8����,ͽz��Nl.�u/z�����,��*�Jh!Ea|]�Jqȁ�3d�}����k$M�$:;TG�[L.�g�R^,F����,V�t^�������$���q?:n��'\�lz>�W8:� a��p~"%��VL�磠x�����5���Ѝ�
)�W?S�s�N#k�ā��4�˘Bzt�RXEz��MW'��p�IW?T�~��H�˔����J��������˸r�ҥփI,"��#��WV��Y�|�@�?��1�����vΦcc&z����EG7��o�ՠ f3ڲ�fi��p��C(�5|O).����/��~O;2g�}U��>�_�Sz�jЁ01KܼM�P�'��B����<���
�,��`��J#�ר~H�:<W��`o���2����)�]���΁�'���5�䄥��ǔ>�����>Lm{i���=M�G�e}@3 h_S=��˥��o��sd�B���}� ���������(Z3�����E(�����7�{��F��O�.�I�"Ů
ٰ*����Fv��?6�|�cQ������!��O����c9^�ա�H�ٮ�D$hҳ?�k!V�2�.��)O�Z���ЯP<xh�D�ͱ��a�"���vG��YǕ�u��/M��,�����V!Q����NP� :����I��$��:6��;��eG�4�j�������Lm�k\�.�E!������������5�H4V��G������X͖���S%7C��V)����P�MøZRK�JsK5's�
�I��C.�ڬ�b*��)�A�ч��}�'"ùj���YV�^���Ѕ�]k�/��s��ۍ(1��E�JH|�A����/@��WU�s6�r���@_>���'�`qq`��J�N`]�ȿ{[eFdG*/�o��G�6�����^c$��ޯtq�$����R�[9����_!�t�G�=��ڿgB�W�ALVV�(�����a�_��PM���$-��b)��X5�z�R����up���i�^V槳�gP��-1�SHM<��e��R��9q���y��KN���ž zļ����ȇ.NO��g��z��I��:���EMx���m��Eu~(	������k
�a�:����<���M�>�p#$/�N�O�)�eh��V��?�j���ٷ����P8�
��س�5���ans]�.�~i.c�߱^O�����/��������%��6I���o�R{�^܋&$���\�֨"��4g�M�z���<8>��ez�w�ؘA�@a�8g�l�tǉE�e����1��A�n���.DP�x��
-m��6#8�OA*_�Ă�#�O���1�l������y))������}��|��r�{���(��ǈ�Q_!9�ޭp3��,@�ӷ�v#�3�C쎌+�HDK�i�Mdhb&� ~�����a����5�)���I\A�43G����5��G=���(�⛑$�Hn�lm��Y+�D�dm�!� �'H��fKL7|���PPK�}���u�?J�܃F%�Y�bY���O�m:f]3Ej��@A�*���^3{���L���)s�֕ώ'/�^�!��]�ծ��Q�G�؅u�{��#!�,��WA���S��
��N2� 1�!��y���dʃ�e"��m�Wa�H��}ǄG=���	L��[�|L��
�B����Yd����n�����`ϩC%Y�_�G)߆[98�W�o?�����Y$�|_�"d�׶������5���DXΉ|a�dE'ܩ�Ϊ�l=����W#Kr�`ϛ�7�o��E4Q ,g���&��TC�B(�x+81|�ǵ�d�!=M��VI����B�^��F�g��&��w6��2�A F�n	W��+�� �v<��׫�cg�L֝$wx���x��L/UG��u������q����b��ӹJ������~dSP�r���e�~Uw(�����H1���=c1_8v����Gw��}�
�>����֞�2��6�y]�JK������]������;U�t�ɻ~��]l�$7�K1����d��V�m��Rm�`��Z����^g��Ɏ�@��:�ޥO���F�k���
�K\+\�B,)�a��Pkk���-����@�Ԕ��[�\Ϙ?�o�#U}���(�pl*�Um����������ME�TN��Hܮwȿ:ɔd��.�G��ㄿ��c�dBsbby�cUy�r�	[��/�~�ven��c>]��&:AG�6O�Z�w��+	��k�܇��	�$'[V�6��ь�eb�����d��;W"{(�PN�1���M��uݷ�'�i��?��J���p��P�r ;�p�]�I���"��Id%�F���5�4�>�2]�A����GN����R#JT5H���&5�'\7�t�z�BO���(p��Q�rp�I�iOt-%YVե����!�V��7]1D���Gl���#Bf�!��|�|�����P���;�:V����\�m8�%�vTp��F��{O6&��b��a�����?Jt�M��-��z9̷�����}[�����Z�و�l�g��T��9���D~e |W,L� �(�� �7����of��#��_�16�D��P�`�R.�"�u����)Y���`w�گĢv�b�w^�aO��~K�Z�T�&N����h�C;�[E�%o0O慺4L���$.�X��Z��\�N=� _��*�6-d�|�0�'��3�$�M�u޹�Se����Q�܅S�����O�w��� �Sm���!2^쁦7L*��:c7lt[���L�)d��!I$0m��C�Ո�0D�rd�p\~W`CD��#wb��܄E��5
d����_U.q�.f���w�n�ޕQ9�`���$Z+��T[n�2��^�.Y+C��:Ϗ-T�#��!�ؼ�J��:$��O�>o<�(�s	Ȋ�:��+��96�b�d�L���t���f��A�j�yH���.|d�l/�lvp�F}9���P��J�-M���}9ѿ��w���&��.v������k�/�
U[h�|_�$h�

�4>���}e%"��H�4 ��r�堝��P�f�2�m��:����5>��tM�[zc����h]��.ɿЫV.�Ȩ����_�R�1���tO>~�l�L-}�)ߋ�&�|F��ܒ�P��u�� b�� �e�5t�� ��U
��U�#��a<�{�4�ӧ�����@�F�iv�R1XuNޮn��A�]��ڿ���l�\p�>c�Vl��]�lbz>̣'z*Ǜ��A���
�m E�C�A��������fM���Ӟ���n��I��Z%̎G��'��U0ͨr�WF��,1���XE#���'#�Pj��Ü���[<ZA'��&
E=l�@ZwKq�������$�W���6��$��w�*�W< �����o��gX`
��f�,<ν�+�Rc����v�٭B$�vx�S?q��`��k�3K��ݘC��꫺.�_��I6k��t�m��rK�:��y�����*|��CjI"�s�|�0>aP�$j�\���O�F���6�y�������h`}�;�������X;�P����m��D�ؐQ�e��ԫS�W�XXT����Ժ	�1~5bY��5���PS[�m�;$�����0Ϭ�W�[�v�\��Q��zz{~I��s��Mq����Oo�E�m}?�u�����i�$(�5Y�@5Eh� F��z��t�0���S�w�Z��te͝(!#�#�ؓ��l��oS8����$���djc�N��!��l�����J��{{�g�N�/;p���E���d�f\����T�� ���7�-j��E�@��z��#��"=��#�s
=`�7��O�d����� �/p1�闧�!�u4�"�r@�����QK����܁дW2���8�L�
���>A�l�V�
-6Up���Ӓ����t|�#�y�Ȳ�T@_���,�Q։�;�Ew�i-'���?E���jTu�J��صܡS���n���˂a����m���I��Y8�m��D�6��O���_6��=̶��d�kX�-�-Xk��f)\��U���T�4T�s5+�7��1����jQ�G��]�?�l�蜾a<�"5} ��̛P>�Оŷ~��/�'�������ɞ�����ٱd���V�I�����F�/y��|�i�uY�=�4�=x5���:�Xƫ-�
b����F�����!�lQ5�(���@8��L)'��Δ`+�qtY2*��3�J��z~��Ie/�pR��	5���7����ЁH����e���zr���oU�t����~GŲ��=H �'�Pdۦ,X��PE�&�^P��5s>p2W	�:��˝��Z�2ױ&�wxb����8�;�+t���l��U�27�v34��������#�/�~;�x�4�bF��H���e�n0��ٓb*�U���$ߠۉ�#�ٳ*�*c��_��N�	��`�2���������N��vM�������(]��P`�A� ��/W*��� NN܃,m+.uπ�!��_(�b�@���o�VbJ��` O�V���Z���z�$AyI������J!^n\���p�kp�#��������r�*����� OP>��!�	&�ǙE*)%H�,�q�3��d �'��w��\
 *ro fħ�!p5�;tЮ���d9i+�w�W��|�2�O(��ST��[J�l������F�uK{Z#X ���vn;j¤��)�ۑ�(���&��J���I�����I��u�K��65���H��n�F熣��T3L����}�Z����˼�o=�Б;�jn+�k����������ElhAgN�U*�\Ǿ��&�N�
ņ��7.ǋ�5��9�g_�\�0��]�#�	<�8 �!6 bÆD�����T��<y���Y���o,�G2�+�0��v"��(�� URK<��Ҳc1��N�`M|yh�cqӴ������ �	�.n�q�却T}�b���<3�C�5��>lcJKע����ې`)��)���G��/x��A�� �X�&!~��.}f��I˴��
�gK���3v`��obTĤ6E��S���bY��L��	,6��=C�%�)5�	l&�ў����?۝���͹0|�ہ�f��q)%���G5���ޘ��k��^79�'�~�~̓�#-�<���CX����(bgY��v������Q�R&���d6mb�]j&�5S,��N5����"(	؀��FB��X�#�1�?{�����^�ޣ�ě4N�8��OE6PA5�����h%�u��������a���w?���TI��@a���6��~��{�u���7/�lTT�ӌ�k�C���9�*<+�e�*�+�u�ϟ�L辰�JR�b���p8%���{gI&��������w�����>ޛ!�82�o�FЁ�슄K�Y�K��ͼ1P{Fg���>�z���Ý��r��U{��]O>^72�vS��؆%(�T�/O�#�bU�]TxJ�ƫW��>��Q��^�ʟ�#��B�޽(r����nֻMP�ס��w	S�Ms�+u~�Q-#?Q/߬���HO9�ɁUZ�4LM\D�>�7���Q2�NSH��%�R��|�չ vJ�
GO�N�_y�sa%B��v�`f�r+�'+<�z-�d�=�����X�z�wA�(����ku�꧝�W�s~���?ˣr�u���$V�q�	�c4M��r�Լd�u��%��O�wD��`�#����f�@��|Z%�'��C���,R	{L2���q��$�f�2�)�Bx��RS�:%��魯�7tCҊ����g���G<���ЂB���Whhz���M���f��E�E��Ө9���h�����x�"1�k�/*�GC0�72Y1 n�[}�Q}�y'���u��9�jb�A�3J$.�i�bq͍7k)_+�C����0��Ƚ�A$">�,uN����o��s��T�6$��/���c�2��}�3�B��&���%�۵�M! �5�fehӝX��ie[�6f���&���%l�<�YçZ���������d��;,�b�Xc��.Lyح��K����XG��S�����\p	5t��J�-���l��q���wF�ͭ�y�3�{x��OPho%N��hq߫���\�?���e�/P8��S��f	�5��[m��1W{�㸗ʗ�"�w�gA�q'Ġ�#C�u]VB����O���� �������`�q���n*�uC����<x��M3mӵ���c#�jhN���7�������ܯz��Ņ�
!Hn�%Mv�V�i�&�p�7-���:s��pV���}>��!Ynz�hSτ뻉,W�8VwN�i������,}��L�R��q\�$Q�- ���m�u5�R�U=[\�ӁM�Q0���@��m]����8����WIR�*�2飩#�a��PgF4F35�*[C�f���0�"옵�����Ht/[A����jo��:��,�Re;����U�ܻ4q��Ӷ��@8ű�
�(h��aQ��$��!�o���C�?;����C �u���N�\/1|������e�Ɣ	�4IA�n2ʡ'�Q7t����nK�r�;�I35l �}�e `T���1�d�
V$��D�#/ۤ�l�yU�UR%��R��	וc瑀�O16U	Qzp�Qv�V�I�2���ȹ�w��o���&����:��t�!�ƾ+���SxlW(aܽ��,'�j=BL`:�6W���C1���n�&��;+`��Kr7Ő���Ğ6t?���Z���̾�ܫ	��Jt�u�ak:�/���$�����q�W���uB���אۍU�Ej�����l��rgKT7���h�#Ҝ@��C�႓�ҿ�c����4�)\;�2�As�Dl
v����5�7	G5G� k�x"�����u{6�r�m�����o��M�<g�/�TǰV��|HQIk�d���h���ŋ7nMJ�5y�	l&
ƣ��;��B�h*�u�h�u�1��t.�D��Y�>�,(fU�}`?��e���v���?z@��]������a93�S+N�M�h+�\�=7�W����Ԡ�ki��vv6.��6� � 2�� ��4E?n������VH���R�,��FV,�}������&PB��{�k}'+�����S-����O�zҿ�)�m\o�������I���°�D"�B&��r��߹?y�w�5-�$K���bQ�]�b���
�ղ��O1"�����7]ʒ@�|շULS�o� $G����`0l��K1J=����(�#�I��Կ� ��W����?|ɳ�/
~�m+���"�]Ys�s%��	�ͮϓ���h�7�b4�ȋ���'�KN��Y�On��Z�O{� 4j�m�&�}����Ë6`ؔ/$�P��{�Mo
��e�O)mT�D�Z�=���`^����b���nk�ۮ���Y���cs�<8�Q;�w걍�c���	&�R����}k����_�3_�˝?������Q6��#�;�mԜ<t�׫�"�7&�x_|0u���%rS����E��� 8�F�q�S;ˠ)Є�~��\��@�P�����X?Z,Ztk4��,��R�]X��i���:l+��u6g�ٲA����V+�E\x]��L7����s�$�y8J��Fpi^h �N������C'wL��P�Sς`F�C���"U�Ng��|����ffUTu�i:DQ@���=��:`$3�	sB�����!���fa����r�:��oz����)#�����K����b��ZP�eB���n,����̈́N�^��n���~��F��'���Ag�9�%Y5�u!Q�/πc=s:�z��2��u``�0�t���j�����ԣh���&��Y�`���w�jo�k�g� h�|6�<����v7E=U>����I5�.a+�^��.gŤ^�"�s�t��n<D�?�J���v�P<;�t�5v�`��GFU��%\F=�4�&�Ь"�����b�&��ٝk�-��v`�a!�(BD=*��;����G�1m=`"�~�$b �!�Vteg�ں7�wly�_bt�f(/ؑ|�x��I
o�f�G7������#��9Hm�	y���m��tN���q�����������^�Img�r>`�ƴb	rp��~O��<4Kܶ�</ΞgܫGS�L���h���C���On�}���c{<��2�=E`D\��o����L�4^J����ap/sh�9���J�f��&�כ�i��R�4�O�9�)����	|��3kpǲ���V�$�Rx��3�����`7��*Aq�nk�I,B@�a����|=���r3�o[<��s�Ů��X�g�G>��"��~���'�;<�c����M��]� ̴O�$�3�s�����v��mH)��k��ɷ�c����@����D=��7� J;{�%��`~¸�R�C/D�_���/ت6���/�yv�W)��>q�R�Ov�Ru2E�܉�C�e]�;
?˝10�uꝋ�(��[�vN)OC�{�!�'�:�6�+�=�q��.6�| 1*a���
(����� 
e8�&Qs�Qp\<�G�wG�'����<�	��"�7Z�A�^x���<�5pw�����i	O��;����p����Gȋ~ҍd�9Fjm<sL�.�L�3k���1&SV��f�t2Ie���9e�N�ۉ�O�I�J��Vܨk���B��j�^`y�w?L)�hA��u�G*ލ]�E��-�B�7���c��U�`6�ap�ެ�����Ì��B;�m,�L�,({��(���ԗ�ӻ��aL&r�4��f����؄�vһ���7k����U9�h�ad��cWZ8���Yߏ�\�'�wrG&S�Ek�F�������~"�U�5y�P��픇P��B8� �]�.�9����ϴ���^��_HT�.�����8�Q�n�e	��Q�0}�6Z-�}6E�T�"E��}�\�9��L���Z	぀��|o`g%Ʊ��Մ��4F�j�Q��Jf��Or ���*��X�,���`"� ���6�)���Lp��(Vdfh'3�X����A|�t�g�L�U)�U����b&"ʌ��!S��CcS�J{�9���bX8p!y�R�-���ԉwe I��*���7�=ޒ{^~ ;=�k �Ct�3�Z^G��-3�Ǉ��L����1i���sx��r7D�ݢ�=�y�hp]!�)�Y�=��w��>�L;�'�y��`+٬u�j�����U~�980IL��������S�aD�����y`�r�jH�	@v� �~#�MW9#iS^ӨЏ0�Y��dd$p��/�5�K�W|v�(����r�^{�3��Te��{�����#B�&�`ֵ��G�E#٩�6��k����&�2�����r�b!F���`JpH�+���M����:�f�V8R�[0��;��x��O�Ʃ�-�B��ߘ����)L\Q��f��T1��JD��^�)r���&��dXq=r�O��ɋ'�a4h����J�R�@�Q�A!�>t(���χ�7�"�_��"m4�a�u�c�i\(�%��ej��\5��:z�Pc�p����> �ʰ��#�%}a:�ώ�P,Y5N�/C�������Y�d��f�`u���iMZu:Y-3D=�9Ʒ����Ό֎�D#�]�;6~0>|�\���e�q�&�4D'�Y�t}B� -�,��m��8���ki0�<�ĺ�6���isj+�r?��y��`���V��( �N��3Jբ�䯵E�GqX╎�\y|���LW����#-f�ۍ~XJ�̐0qe$��ó�c�Y�
I�^׍r��H�$Ypi�QV��B~�� u�G@'�^;��S髝f�a��BI� ���۴ǆT�!��p��Qh�]�;���-S�,,�[IH8�[?�Gg����C;�
�*�`9Z��5�PhJ�ދ���Jt0>q7h|[�FY����JQ�F�[ӗ�9�G��V���g�k�65-�};)�b�i_ˏ�߱G�pDi�bs�w'������i��adqW_�5���q�Qkh��ʴh��[�2(�J"lR��e�����3O��$��U%k�C�'�豛���r�K��������8�"���Q�+p����x� �sy_p@%���� 碢��N���O�C��Da�H�)��P��n�g�+�ʯӲ\��B&���3���ȵG�L�r����ޱl�bV�h��䨞�'3���n�~x��'�[8�l��/�����k;����f؋��c6�«�FX��*$B��W&�R�v_"�1>y�K꽲��u#aK�'Z����*�Vϭ%A{������I^y�GY"��K�v*�Gaf}'��ǰd�/� ��#١@�x��	+ɖ�2���*?J �usĴyQ�ʆ�� �O�b?�ө~ƣ��CV7���}wE 32$����C54��YP؄VN	�*�ݵ��I�����.G�
����z�(os!������UHVN��ӭI�  �pP�\! }O̓���[�Px�)�|�^����/,v'&q�.���������-G#�A�`�+�@���_��-g��_�GN1�du�yu��h�
��gμ�f�UT|l�E���?�t?�ҭ ���tWrJ2��ۋ���QGn���g#ӧ�;��>m���)�-n1|��_��N����s��ݱ�#���Ħ�M�pl Á���u�ck��]�&Җ�8/�(#���x	�1����ӼD����)�x5����T�#�GbP$�1��;D�����m&��{�Vb�.2����e�G��#-��$���x���td��^��W"�$jJj�����*%�������?�`���ī�5��p�xΟG�j@�nÏ�4⋡>`�V�
嬁2��E{�y�J�r �{���dG?���Zy
Nf���D�<���g�C�^��zG���B��.�
:�z_~�M
! D�iBT(r�p5��$�ST=F"2�8�Γ�	��c��-�(3f�jh�#�[=�.�вܤ�P2��'�e×�V@�����UD"ny��G꧋?���B�A�M"������_��J
��7 b�mA�WB-��?�K�N�6��:Lu)>�4,�1^�3-J_�)И4��4BY�l��*׫����������J��
#p��!��Lc�C]�(��4J����f����;��o����_3�լ�`[�w�5h޾z���b����`��5��^iB,0�@?C��˒�^`�{*�Ӭ4���gI����60u��ؿk�/���ִ�i�'I��|^�  ����O翎Ɣ'�N��"���725�/��ɀ�_ � ��򖡮3U��Ui�������cr��*c*�q��o\L�1>Nˉ� �NN��6,�g���!֒��nQ��Y{����!��Y��向�Ql��Cq����Ws�ury$*�bȞ3׳���