��/  t3�k��Z���E=@�D���*8|UNu��*j���*S���`�2U�Q��b�x���W*��-���]�0p� j��b����i8��Z�<(��žz�#ٔ�в�v)/�v������E�b���F�;�^�xK"񰾩[���dI�hz��� �%܋�s^��<�J���
U%�F�}�(����pE���]������W
��/]��ҭ��oE�F{��\�b�ų`@�P��C�� _m�!ud���/�ݢ�
�7޻.����P4��s�i�\>`�@�u)���f��2J����"���Ca����6t�)xG���L�-����l�V��)�2�-����\(@q��V����C�>8��#w`g	��|�G��/;�&����y��J{@�v�K�+��i�ٞWI�|98�U���l�Y�C"��LqyP��U�z|�Uo��+���K�0��\��� �:�����Q_����G��}թ����2����O���t}Q��$������9o$�v#?S��{������u�#O�y�L�iZG2��u���P�W<eK���6oG�h���G���쒹��>��k��J�IR��JR����K1�U=H"+���/^T�/�t=��OLt��1��3:o�ĠU��z� s�9Vz�C�AuCج���}�w8����JrO�G���N����a)& u'y�^G�F���5Ϻi�H�D+0L2�ܱk|W�{	�h�Wl�<�[I�&wS-0w��;�_��yՑ�M��R�s�]��ajQ���B���8�A��\�ȉj2L�3���$j����L�����Pq�3�	�6�nr��V5"eV��*O�h�RT6����^G58Zraj��w��<Y�"��]��,,�Ui�~����s��Y�����ϓH�v�E����~��ܻE2C��[*}{W�C��4@T���Kt�%��ӹ�W�S[��^�̥(�bMQ�j�(t��j9W|j���"���<�����'�!JW���xXE4� �L5ɖU����q�g̽��tGӎ�������E�����HL�'En��f����DDE|c�~�]1|�_O:�'N�|�=���.��5��~�D_N휊2�����r;}װ��?�P�� ����ј��B5����+����2f��5��|��3����������e	<�%o�Y��ʌ�Y�w��T��A&+#I�0� ����\�a~���R����������ѻ��a�TP�Q�p�P��LY���vċ�8t���a�5����i����F����	�JM����c��,Fꐸ�j *3OvW�(k�	̦� �z��>���\���D�Vo������@{���v�l���@���\�Yu4E��Ll�7�\�W�Qf�X$�6L�b߸��;�69C��c`�l�+�8����O�q���&m_�ev�<��P ˷�֥;�~vK��FaA�'%��&m&�F#��?��%Rdu�;y���a�����+	�������[�?߹j�Oq^|��m��/Y��M�F�G�}�����g�-v-�KgX_�v�Z]�y��[�ű���f��C���i:L����a��g�C���"!�?�xAN|D�AT��E�G ��!��Ԍxb"i��tT��Q�liUD���wz�N����6�A�6���0q���À7��� �=]'�Ou��Ch���'� �b��?����ӓI�����EV҉�]�`��״(O�:�x��i%��rm&����P�gN�@ʒ/0^搏��%<���a��
��(bD��N(�m7�6qK��;$��.2	�ah�'�3�~J�
z %��-��N?�d���f��h*gk�����m���H�SD��c���'�JRo�v�:��vZ��3$V]��je Ž$� ŴE5NH����m�����`��ޅP��|�3[�_a�p�^ۃ��o��D�4��w�-��R�V����&!E��T7�Q�y(�[ڤ��ܵ!��J��?�jjW�30��zVV��@[�Α%�ɠ��"-1�:Zɍ�Ү�����4�-l�����n@�v5��-w��5]���<�(��X��]d���wL���&����b�%⪎�˞�
��A	%T�||���R����m��ԋKaU7�_t0��c��k�i�Zv��E�&Ѡ�j�=�V�r���ٟ{7�qv)_��5�N5�aUJ)ʷ���ul4�@o�;i��R`���b��&g���=^�O�{���b�3. ��o�����5�r���l���8R?�?����'���{�}nGl	;�\� AaȢ���t�.7�-"d>h���@h�}�],���|d�})��N�?�k� ȆV��X��&�4��)���̨_u�fΉ5<�1}��Z�hy
���ԣ3&��� ��5ǅd��N�0J<��+��ن���%D`���{�I|��2~
�eXȤ܇�mq��IZ���e�C�x$1&�'��$M׳ ,��?܉Y+	T����Z>i��M�C�<�OZ�/��+�{9�@?�����X��a�o�a��V�&���G�0�zv7�!��X��⏜vR��v:͡��罎t�㼊T�rT�5DC�J�r��(���G���]l]l��C��)�et�~��M~$�R�^H�4sz�Ư��l<�b�h1�"q��P�&�L���"N�8�,��9o�#Kߺ� �Z�$j�����{!	f�
�h��^\	��q��t#��iNJH��ݸ��goY?��M�W���u}\�U�;�&�%���&���M�*�aតz);jV��̈�-Qwb$L�W4�{���r���\��;�y��:���(��6O�a+���L��p�]0"����Ғ(� D�b>�ov�w�=��=�����4�0�鏋��t�*9k;"C:����e#�0�H��mƺM~�z���,ef���p_%/e-����*{O�o�*6��c���9���1[��]qx$���֕��i�a�dr��M�­�B:
�M�%���:�J�rK�&D�{��2������l���_,�*c�
i��o��H�0_��^V/��J��+�#��P�[M�I����)��̒�� �Y�"����1��$�_[�a�U��KQ:d}��1��/��q-_�1�EP������k;%"d�y����/}]`hZojjA�먟�➰�`���-hT6>�h�Q�u�JX�<��$SH�d�^kxg�dg����rԠ˟���F���Q#���&�`���afC���!�X��V鰓��]�^�+��OY0������.�h2��uϬ�=��kk���Sܮ_���P�X��`����1utZ�C��!уz��;��!��!��� �����K |e��F>\QC)����*�v��Hiϸ#`z������jdF�T�����*,�5sx��4,c�p�,ͺ�B���`N�6�f"L����|���f1G䮪|r�z[��h],VP%�Ƀ/��_���I�l�í�����'�靑�olqu�tQm9>���l�v:�6UC������}�94�e~a��o�h�.g�-����r�j55�H��<���9<l� � �e���l.d�c�U������`=��]���훋���QQ�A���H��2�)��о � (��kO{�F�ij8�E�P!�
�	saD��4� ��_v�\5�-@Q�Ϧ��bX�b0k�0Ș:=M�*❌�U�C�m��L��܀!O�-f�M�p��A�#�������㋚�r���b� ���+��S��Wk(�+��8O���zW���U� A]1Q��]_4j�X9��;_F�?M9	47�8�q5�#b���>�lWl|9!у��]I���_P,&RF���h��k�lq�ُ��o�P2��1��pY�f��eB���2�|�ir�So��@)zժ���*���4)�Ū�ه�%Ɖ���J��]z&:S^ʒ�6�'�h��^��*���ׂQ���=i�~�Ƃ�)6w���G�< KB�wT����՜�N�|]���,2�7�*�K���<	�!�f�*���T@@fw<�C�'��[��ۺ��I��Q��<i��5��se��+u=�(�]+N3��ο��:��^;��$,.�I`SI�XL�ꫲ�����Q��	�1]�S^0<a;7��k�Y�����	Aڑ}�	X<4��r��>��g�Zȧ�@�8+�Q� �3��;L5��f��f|2��%j
�PT��m��vl�M�`Zn����7>�Y���pNܷbm)�9��δ�]���E���Lf��%�\����� ��p2�z�����m��B� �$M��M_%WY*i��W�n� �޵�Ⱥ�:��.h��z|��fU�'�0M���S7>T+�6ބ�(�?xn�̡��w"4�{��[B��\�S�M/3�>|��׼s����1_Q�9��L�*������M���.�S%�.Vb��`xiŞݪ7:���Yޫx/U���q�y��`{Xo�Y�s���%�cT������ti�_���>�a��*DAA`����E_0��"'Դ젰rSG*:�?�qJ�(��ӭ3�9ct��Z�oĽ!���k�䄧|��`����.N~j�[�
�%���(�Z>W}�0���%��l�[9���n=�'�|����g叮 ՠ�z�������M�?\r�����L���9�>���x��OUv�sR��O�H����D6�����@��Gˬ �u׬.�����+%Q\���'������U0
�3)M�I0�U�k�$č/ف��HaK�v�4r?�K���X��z��I�;��]c��{�rv���:��qꃐ���њ�q�x��z�Mܾ�H�8ԉx�!^'9*�s-��AY`=��� ��a�)�ӦU�I;4u�@�n�sH��>�N�I����(ID�� �
G��E2Q���>G�����!�ʼ���	͝��V�#I*�#����o��H>ܰ��2�{�mC6��n�q�������{</-�Dװ��a����蹶�a�pG�S$�
ig�bf�Zdk��y����wy��|Yȹz~�f��g><����Fy�{i�PN��f�t�ml&-���4���=�	Ɓz��X`,��� �V2��:U�E���")�ѓw�/�U�Z���K�/A�ʏ��;$�8��E�e=qf_T=�%a��P��UP� �jڦ�/��<�~��ש	˸�S����Wn��r:*v*��Zk�(��!���r�G�j)oψ�<AUN��I"J�߫r��q!�y1�2 ��\��L([�ZŤd���=Une9Q>c�Adk�`HՍ���l.Nyܚ��:c:��i��X�3c�B���|�������"AB��Lx1Orz�����t۵���8��D;�n�yF��P�l�Ms#x�1"����f����Y0�s*E�z����>�g>��;1���.�Mt;	����.�E�������wo���>��CF6ٻ���YN�,��BXWP"�7J�fv�>����-\�P�u|�Qb����_2�ȄVj�ol9?�6�Ż�KH@9u���]�F�R��?���%��Tg����%�`�����U2��p҇<m>BѮ���W�u�(�Z��93��d���1sf�$�Gl�����%)�=b��mJD?��$��(�!TQ����O���l]��$P=`�I���Vd�i�2���!}S^3���C�z[s�
��_���fq5�M����7��-y+���O[p6eߙ+�2�	��Ù�×hb�<�t����h�{i%5XQ��WK���M����[<*Ú9��3#]Ժ�\�I�sk�e��HA��W�saJ�[2���6mXa�{/K��s�Tʉ����ߣM�?�X�r�W��g�v��
<g�c�L��{=�F��cR��Z���R/����|�.O<,T
P�"iX���_9��)o���`sr�ǽ3� -x�ԃw<[
X���^FPV�:�ܫjv^ 	�6�\V�J�<f��S�R�f�������A-�����c��Dō8�PK�5ځ�G��e8*.7ժ�hȟ1��"�[aR+����Ы����n\;A��>���Q�b �:�]Sjb�#��0X{n����#U[�Bc���:փ����ǖ+m�e��W;r���|�(��ٍ�Kw�ھ	�KP��Rūi�Ҝ���n�c���XbЯZ��[�p�a8�Dp������ۡ�x�ax�!P]~F�2�w�0���� ��bہ.������˽u�%��]�5 �'�B���Vxۻ��+]�i2�K)����l�eo9l���տ��m�Q;S�'ų_~�٬57�?�>�hYj�@�*��cwv#�������]v�K=09�T�/��q9/Ha̭���mJ�k�KNwEYT-0�̓@���ZzR�R�l딈��|����]�Z�V��ȯ�`��00�$3WkRz��'��Œ?Ǳx��[�6}i�4��õ��E��+�_�$�(Le��]V�i^2�Ve��r,���@���q =U���
Q����%5�q���Td��D�TG���<����C��hLϧ� �����6�)�9I7Ckz���	z,��IP f��F�|�f=�H[��0D���0���Eoߗ�qEu�� )r%��hFq^�w:�^i��=�uP�!8��~��5�jMO�R>���m(|�ҵ��B7#8�K��d��d��`À`�!{&�Gi�w=ԫX�O5��	kX,�^��:lJ�[�.1��#E���l�W�k���r¢F&���e��kˎ�A]�v��w(� /�~��>@˛��&8όju{�j��i��yΉ 5K���)��,��f�@k��d���Psx��6[����h�����i�� �;��>3�y�4��:1AY��F&������yo?I.g�2��;�E��Y� � ��G"���(<����Lq<V������Ǻ�-t����v1
l�׾�����jZB�cp�EZ��<�j��̹���p����o��m)e{fԢ��[sӟ��s�(2Z�TB1��0nFa�(��k��ȶ>T�Wj�" 1� o�Z;08npw^�&<��u�t�&�
�&�$D9ݫMb</1�2c����Khf�1≏�.����:�ڟ�)I�A�ͳ�4|i^4�uĩ�!�vm�y�A�m]��&>�b���(VU�G^���5>
�UϽ�c�v�]}�؊�7�"!û�<����$Q$>�Q�0�P�އͫ�gu�����٘a����L&v�wl�p,7S)4�S,{��+���Yu�K�[!�o��`��<���7�Q�?]\���ܱtJ;��xn��u�_ú�qCw�%=M0W�����q��cc��*�`��=T^`Z\�x�i?,�R�CG;��#�As�����(�Y]��Aۡ�}-�������N�/�>�.�D�z7�.�\K�J�ݩ���{���ɻ`y��H�6S]E���ZJ8�~��}M�(� ��~������Y���$�"($��h(o�׈��\dx�f��R�: ����f����G
�l��8ǐ	x�����z��r��\�7k#u}}��c.�����c�U�*9Q��z�ή�"5��֩F�@K��$��C]�YH��i�fV���C}n�e�o�.f~�����Z�%l%�q����v$��.���T�-�Q�xKr�1�ԞB�o�`5Q�S?�[�s��|0N��n��Ggڞ��mR�$z"K�N?��{	�6>�L �'�	ֲ:�b�C@x`��gn�q���εh�3g�"˰U�>$^X�>랒b��2�EQ��:=Ŏۃ�g�	���R���f<�\uXP��eڄ�B9^�#�W	hS��3f�)6��`$wF����>���p�.��"*�|@ϴApk-]��7f�#�A���x����]�_^���@�6s��d���_'���UC�Opd�ջ��!�9������x�F��i�ť2)a�uMH��N����h�bdը�-S}�� �?�庅�U/�?���|�C��luW�_:�,;���\>�Y�
`\1]Cw��!,Fsڔ"��M�K��ҳ����Y���I���UN� �m�����V�;ɓ�E���ʴ3 ��'�M���Q�\`� ['Ń7�u:��-vNL)L�o{��'��O�L�ܯ�s�;b�.�ā$��'� �xXz 1
���9�.�k�{ASj��R
�Qkkf�<��t�3oSk��Tm�3g�hS�Yg�t���%�צL� *Vܓ� �*�E�����O�8��Lܒ|��ŐH;z �|��r���x���-�H�����7�7@�ٳ�ނ�FM�Pv�yU_*�9�9��=Lu�_�E@]Wؒa��ASg?@6��)�('�r��F�u�����.Fif.�v�����i��\�
�N��a�'���"I����밡�A�x@*��Q�X~e���""�+�i���t��<��.�AT��"��>���׈ښ�b����_Xa��7�E�Ƶ�k���ed`]�ey�C�����q�5I�f3�׏�U`���$@���u���܁��.�!>mw.9�^|�'֯Q�zU$��.@}��^G�+D�l�$��I�����5O��ܲ�ݍ��2K����瘼�cQAC;�P�:БC�ƍ�K���hM��l�V�_���)��I��b�C�^h^�j֖�݊�Qm�mL�4�ޫ>J�!0��Z����Ig����n�v��J*�f��zEi��M:%>I�P�Y���N��{i��d�xJ!2����~fn&!A��@;�3��'�HtF4��m��:��s�ƭ��R��ԟ�%�ˑ��!��%wג���³~��Bm�p麇��7��Hj�/������shu��a�ܧշ�*&�|]���{4�6ؘX��M���NA����d�p�\qD0�w|���q���7
�Q�-�l ]��$�MJ%�u&����P��	V_�,�;�1���5�b�1�Os�3�]�J��-��+Mz��{�G�W�Ĕ�d���S`�c<�����z�}����}��*��K�L¨�:�b�3p�8z�3���6�g�)h1n���[ϲ֎˸m4�`J�h�I�*'u�T9��:��>��!���GCq�kJ��E��/�-��|ډ��F�A ��2E�L�5��5�"߁�g�-r��'�nc�k>�	�θ@��DM�"W��~�g_H$��q��0s��P_G��xכ�=��
q��Q�r���sHf�����c�����Wڇ?^f��@��}�\1���7�_�W8��0���Q��s���t?U�I�?�;�4�������!�9y��`/>�+'1POL�d8v����z��5�GV�=CǊ��Q0��,��J����e>���o,O_R}���LPY9
�s�{��ā���	�,��#�$y7���_"(_3�=y<k^:b�r�
Ȉ)�j�r� �6�ts��4��dy\��<ˎD�tN��x���!��Ε�_�����
V�q�`�X'��x:�6_ sX]U6O�[M�w	��f��iPd"S�Kz��&rƑ0s��M��Omn�����.�{ר�'��Ԫ�oT�["X��{���0}��j8r�M�߭ cJ���>|����w|>�*�$�4U�}��c<�l��\:�7D8���R��Z�uH���_B��C�[ ^�n4] ��[8��M���K[g�#sF�Q����|�@o{I� *Y��7:�2��L�%�$�sN2������߻��MߏVtQ��Z���vǸ�q/۪6�MK����� _O��~�N(�&F�nl��8j�����ᥒ
)�=Dc������~�7��ܣ���ƝKz"����<�#�]ao�i��'iJ.���k�`��a1��8^�S�({������ Y�Ep>o����L�t?ux�\�!R5���G�����2�u )�1>x�-���3T��m�>_!|)鹾���Z��xe���j�,������\Qp��x@t�\���X�����o,�'z:g�e��;y_�ɍ7�^"ׅ4{o��T>،��r����fL^�y�+v'C�������j4c&��_s6���x4�'��@��}�*��+�,��.9�|�A��V���V|�hlu��PWwN3�/�v�9V�`?I�Τ�M:iXY��v�se��y��^�,�Y��D�KY�i�2z�Jt������~BG�*(�hO+��i�蘆7�״�;���gg����R��t��#�0����.�e'��8��C����#�}M�ң������=5	�[!,���d��HjQ4N[]����t�ĭ��a:AqէD`�ĭf�g<���<[f>|ĸgF(��O�uC��5f4�2Z��n��d�����p�ݎ���Y��ѹ����V��o�cK�Ow4�;��>b��4����$�*��7?�ʽX����y�<d��=�w��H\�aiNa�r ��,p���
�ܱ�t�,q�¼>(1�D A�����ǌ9\�B�w2�v�$H$G�w����R�Nk��v����p,z���v�vޫ�h��p�ː3{0J���
���",��C�!�V#s��8�&9�xB+B��Y�"��za���h�"L��52	�Ĉu��}�Ui7�`Ӫڧ����6�NŔ`���`w�R�	/�4��z�Z�ͷX�/�4Ө�����֟���2��QT�K���� ��N��:ܦ:� ���6!I)GG��OOB�q�K�;0'��^:C`���(��JD����i�]� N>i�U�ħd��4�H��v�~Աi���_���U��m�ŧ�3�͂P8��V���A�p����-���n���@�I𐛦�{�#�R�S#,!�ۼ���p�A�EBY&y[��! �t����W��FZ�l�cW}3>��C�E��[��\MB�7�7��:���1���I�N?�O;�߁⼊#�.���\�u��(,5���0�!����n�,[ڜ�n�lh��0�(�(N��R<Vp��|�&��s�N���GD�;���մw���Q��u 8�6b���n��e��)5|[���r7����������_e�V!�N$/�M���(�����X �Ie����׮&�/�K�,y��Ф%e�F����Ώ�I����aL���7�N���l_��b�9�զ�	k���]��6�a��
��1b߾�nup�by�1��-��l�fY\�&Fc|����ɾ��L6��H���J��߾��\��y5�W
�WN`������$V�4n6Ɇ���}c���z����^'Ӡ'�DS�<�ʰ��ˤ,�����B�k�X�=��ã��J2��u�S�y���;�w���U�!/����)tL�J���(�t�T����y��#۵�m�b�����D���~��:�%Ή�H�k)��c��������G,7s��+���ƹ�(���+M�X	���#km
.�irM�0�a��`���>0�*�7��3�S��rSƌ�<6�8Зy��b|7���Od�2�k�����#Z+[�gv�5o���	s���
vfd)E��Oė�N�{�ےa��9RJ�*�B��3�S6-2��烓۶ת��N�|r�bH�l�p�5)���Ŭ�nC~�M��Z_܎Nr�=�\[gJTiYr��\��Q�x���nb|K�(D�2b�pin�ȉW���)t����P�x�(�6.Z�9�5Q��v��
���G�|�)w���799Gy��QWS��������r��[�1@:�*^��
��	��R�rXP3�*�v�~�a�����E�;Q�T�ò+}��HK�
�~�@1�u#�I%B�f�9jR����:+��W�2����)r��3F�[�0�w����i��G](�w�8H�h�%�����==�b=X�vqB����5Q����`	>|W.�%��4���j�|�nv]g=��]V٠��F���l��	G�����>�M��ÎV��*�T]� :4Tut�ذ������1��c��I=H�38��M������x_�	�:9C��v��Rܳ.k��$�]A�ݍ��;��79��D�+(6�+�`�r�N�{�l�J�U����Ӗ�+���_Ų3BY�7�e�8~Z���ΰp�M���/Df�mT��A�c�w:!�~	tv��8�]� �?�t\�g��b��p���io�n��-���y��޵3G��Lܦ��g����"X�"jX9��e�0�mq�F�V��򏎹S��wx9Gk�>�`0f-���FFa\h���A��{����L��>���\I�u,R~��J,2zZ�&n;��3��ܑ��3�07�y���uIˎ~^ X ݽ&��5��Q���S�u8:H�e�Pm�fTI���\5P�p$Ȧ1nĠ�����3^�0M��-���[F��-���yW1��ֳ���Y�^j@��L���h4�J��'謣%<�H���lR\e�S�s��9�r9������	|�L�4�e����>��t;8����r����pZ���|�̳�C⡧Ճ�M�Dl0�T2+$�U�?̶!5(2�J�-c&*�ut���COh����:q}���)9%׭�A!�K<�����!*��5�c^R��ň��O,����Ǽ������F5����x`�vӹ�%8&	��,�(��}Ǥ�=)�������բ�pLp��T|�tu����+����%��4rge�+RU�,����oK��
���`�򕙸zI�m����a���d���l�|��Jۭ*h.��*�9��0�$�Ve�m�[N%�FԺ=�N`�b׬�C1�����-_O����-� N��"`�qt#�p��ZG6��ʉ��@��u��=��_c�=���>@;O�������aQ���a���nT0����[�H+�'�C��imR��'{�/C��k�X*<���b��9�
85����XЪ�}��$��X݀�0�bs�I䲨�VTF��6�|ͤ���3�,]�+��(1ܤ�����r��N ��?��L�Yl��۔&��˷��2��li��0S�2&K`)+g�q��O��LDYg����u���̈́N������4a{�XH��'�������#FrF�α�>���˻��!��b��N��i�k�t�V�&����m \i��a�����p{[b�v�
��ǈ�j+�*˲�'���4�c7�޲ug���tO�����Z?�pLi6[�xaq�MW�y�f7��{�y�TU	���&�G����������E�e[�v��lYd��حs�T���	��d��M��@���̷(}#yՂ���sJ�v�M$���W7�4��3�n�}6H�����Հ�Z���� �������Z5��\r����k0W��K�j�.��SgP1��S���
�������ju��B5�����%�˛�X	ؤ�4ݩ*Y��)��~=�^x/o]\60꠱O��H��"���z�Q�ʏA�CZ�{�k~��92�bs������>�@?��r��x�フ`2z���K.Q��H6c_��+"��x�&8W���*�6I���+��I�?���L����� s'ʗ��e֨w���t������7J�u�`$o�m���~�U�aa�e� �uRolP��(P����$�r�IkH�R,�����Z�(�8C�\�C��Ce���w��'P8w�&N�8����Ά���n�u.x�����
\t���;�ļ~֑s`yy����~DȐ��:�`�ĭ�k�\{sZ��K"��0�@����2��>�������/�Dj}ՎCj�S������d�1���8��!�@��r���������E�_2{e��\�^�W����K u&��Q�c��E?�Q���Y�s�uE�o�/��;��
IM�(yDz
���Ѯ������c�7q��}���|�Z2<�2�Ϊ�%���t�=�����!�[�c��x�ĩ�!���z~�es��;B	l��ʓ��<ss�R�{��W�F�S��������ۥ]�=�U�'��=:�֪Y���.�^�#�]���6<�M��NRϏ�V�(���逰H�h�м�^��V���!���nF��T�)dȕ�}�o�yF9�*�4�}�s5��\*�~�T݇�jk($�:`2���L�p)*�ZV	�Qt#�]�A��R��Ho�m�3~���@J)�v��D��)#}?�w��YaьfE�/�]7��\>��D��l�S�'�*  q`T{_&(]�b������G���w�c�����@�z�
�z�p�-4�l%��'�H�8`���ϐ��H�-�(��:���$�˯1�x���z29��yDs��%/��s������UX4�3t����A%
d� V�O���K}S�H�x1�c��d�|P��߾QW�'ڄ���+z�]�\�1&�R�yC� ��m2C@��v����6pO�O�(�MX�
̪PN���]�G�6Xɪ&O]ecR!�%�}�K㇧|G��7C�l!�~�h2L�?Șt�Gȁ�K�������on��c�2��Ա:Z�'���dP̤�H��4r��+Pa;�`��^�P����K֥D)=*�S��P˵	y^ݱ�A��X���S��D4^mk�D(��$�����7�~"8�����_�Iģ��@�lߓ�1=�k1��M��@�r>}��?,Qհ��bs����r}J�`��~�v/I�ݢ��zԦv2�N�W��>�6�к��l�Q0�n}��=��,�$-�OP"ǯ"N�*$Y
Ql�[���2�QĿ845�����<n��e�o�%��m"i2�p��.�n�8��h�{�%0�u��$��Ʀ!A��;���q��%ei���\i��i���	�}\�:�!�GL��I[�I��%XF���e�)�f��x/�'���va-ny��L<P�6��?��L�j��F�(0-��l#k~�R�\�c�c0Q]���ħ�\��tG���+�6N�z
8�؏� �ק��b0�F���$�a�%f��m*Dq�R�I�TQ��wE��Z��V�9�\�D��.kI�:���
,�$b^�f,�m�����u����M)Y`O�����a߮9�b���Iݐ,�^G��?g6)Zz�.}���_��U{|�R��7_��[a5GqK+����ir�c�[�,z�K4Tf�N��K6r�刄��B�z?�v�k�������i߹���`\G1�0]����M�s��v�E(k8Y��X
C!`AgG�?�֟ݎ�E��!�z�eW�!��~F;*x��&������)Z��!��QD��}w�{�K�Zx&e�i�o�Ab�v��O���^�/u������"v8��jP��&���z�����țڈ�%��z�[ۤ�\/�s�7 #L�0e%O*�})V��#Q�9�G��?�˫��i�5J��p�ͿnVU�yC@^逹?�y�B�L����@u?��b}�{`����&4G��
�����ddv�+J����!�0�r��(�G�c��%�����i)IX����µ}�����4I��F�"�0�I���m|`��o�X��d����y��̻��"��1�-��1��#���;%M�k�+�q����c�2/��w5]�e^ۧ$����C��ai0��<H�V���>��	�ca����LT�����v 3oᶆWa����]箯{�0���v��BJi�rf��/D\H:fJ���F�D�t��u�4y ˜�+�u$޳��#�
��ut��|h	���	��sRKÿZV�ا1VAk�(���M���&\�>��)zi1/T޽랜���4�f3W��|�S�h��;�A!n�kU�K@ʻ<9�эeh8(5ځ�6��ދ��["���7$��-��8�m?PR(�T���:���:��}�bg��}��$�(�7�$�>�d37�?����{��ն����E�����;����og��ǵ��2�f�hM0Q�gF�d:d=ԣ���@`퟾��9%��a���J��GD�[ptW��ܝ �/'U�2/ׁV6@@w��p5�����=����sa!���WH!�<�i<�I�CZq�^CQ�9������Fڷ������ ̺`�~������I)D"�zΑ$�#Ptq����W���E�\b�=���dcf��Ј�C�٘��搘�o�nBJ�rx]�_���c �><��fW����;x��m	�x6��Y�#,  ���D�ܷw��%�d�HݧP��9����!���s�Ze]~�V0�djϞ	]�t���g0*���� ��[Q⿛{�����D ϖ�S�|�[@��{}aX��u+�؈K�j�9������%ҵϾ�≔HP�_�}ْ�$�v*y�S�*�C��*�V����w�*c��Ĳ��X/�R~@Ẁ����^�ִt�'�=0e�T�V~su|Ìk�M�@�o%B���G�£}�MI�H_A&�h�z����`+���:tE
�]�C0��?�
�=$9�?���B�9B�iۅ�8ο�(r�i=V�`CGJ�CD�ctğC>���#d�?��N�A�;���hKht;0�Cd;��<	倜��x�)���=`B��z���^V���xg<t�~��%?qA�A����
d���w������r����|�t��Z���Z���Q�x���}�?�m~��8��&�v�����0�=��^KrLK�i�1sAJ�08I�����8����kj�WM<"�58yJ�ণ�8`�h�~"���9�y=�]G���[o\�I�ɘTǮ��J�p�dk���*<-�-�@�dnD�����Fz��1'��xe40�A�L[X��e�T��c3�������d���&�.�	��'�.�~k2�r�`�~�.)� ��[d�s��t�p��m��-�l�������d��kh���O}*�f�4����v��6i���jϕ� ����}�ܚ��r����ժ��<	��g 1.B�H��u��1HC��m :	hYu��
��D�L���.�n�P�H5�߲dRW���KfR�B!����3z���z72��Uq�fG�Z�9�Y�i��=l�wQ�����Bt���!�}Ȼ2���������DY�f�T�!��0����\�$Jq��c��tޤKįg]�.��n�rq;��x�Fss�ZL4Q����s�mΫ��l�!�����lJ]jO�'���_����$��A�����n#b��ǎ7��y[�`��ڐ�I�<+76O� s�Kq����_�4��CKȣ��ms�DoG��M���-�@��P��#����I�<qE���c�}���(�[�������(�b��D�*�5٢!S=&H��+=v������6ËI^�屲 l��F �-ѝjC ���AB +�e�V]��O�8O߭ZfQ����D�=��a�@���Z�:�v��u�c�~A��`�lsv�ﾲ?�b�YĚ�ɰ�z�˔g�sF1��m����PK�#n�z�Z
0��槑M�����Wv$vzb��E�2!y������&j�g�:�.���8?a3RD��
�ɿ��_ 넜@��sZe�_��?�ά�E����Ð�����Ez����=�D�u'����.s�N�yU!oy��{č�xy��P�l�s*�[�
U�Kx�E��ٓ-���]����Ɣ��ka�����Z|�~�>6�����O����}|��s�����^��M���q�>����9�D�ćg%W�� (�#fg_BQ���Eu���������bX�۹^R�Ł55u��p*�\p}�f�����ON!�U���#�·����Mᖿz���A�[�1ASnU���@�O3z���xL3e� +��x&����<�����s,�q>Ί�Z���g�D�=�s��Zì�=a��p�<,X���]�,^wuu$k���{]��%��ΰP���r'���.Y.���\��,Lxu��bz����� ��5h=�o�ܼ�e�H>s��d�K��2g���;d��j3S�� &ƢW.�;�n^y���(.�U�\����ޢ*A沔�hd����b'q�!�Bõ��݋�=.�6[�}��If�.Y�8\`�{]1��.텰�ϋT(����X+������[2q��d�փ�N�~�H���ui�p�VALz����5.�G9n@,S��È%cv�g�)ϷF-[腿3�������n�q�I���߳!c�|CT�[�C��	�v9�zp��Y�]!��TTROc��.ʮ��i?�sn	R�+� RZ.�KoقT7�d׼�C�W�A��8Z��T �n�/��o�h�E�Hih�Q��F��o�\Y2��:�����y�$E=I|L=j��Ě�a�@�O�R	,连hr?�4������p��2�D��f��>��T�+�T�Q�&�����qF���,���b��z�����5���32��X�{;�z�25T�7�� Xl_̩���Q{������#�e�\�#_�e-�Z����p��հ�Ꮿ���$;�H����X(F�4�azߵC��A�<�RU%ZH-�t"i�����m�Nm��z���e,��7�M��d5��]�i#����؜��Y�2g�- {��#���^��VV0��}mL���Iw%�l�rn\��7�8��YPD*"Y7%}��_;t~,5�:�8������#m�yBpV��n�*h|�b�j�Ǔ�S���K[�+|�Xp>��?�����;�7���z���n�^��F�����!�Zi��.�W�����X�r� Gh���$m�~DYt�j���;��f6o��B�Z���zi�p�Z@ϳ�bo�r�¬<^u��.�3us�k�=����"b�+� ��Ķ 0U�MԆ��2�@�ش�Kk��?vV����|]�r��������$n�0�Ĵ0v�7����#��t�-�ԧՓf�����s�%'�H���1�����ߊ��j]�P=3@S��v�� �a�K�JH�����l8��h]їN�����i�����r�&�	�������g��h��7�k�+�n�,����C}f��M�;U���-��w��o��3�x��gX���Mx��e���7�)��r�M�V�ɟ|��[���MB��a�1���gO̝��^�.H`Ǭ?MBj}��"��!������X0�޺�����k �-�3������`�.�U�^8��^s���ph�+��_�����(1�S�ɢ.�i���!��Q#n���J�P-C���f%��}��M������BF;U�DY��8 ~O���#�*EZp�oW�j��jO̄M��@�ޛ�{�ENp"³�Ĳ�CZ��)�첷�&Q��~�x*Ń�D����zI7��{���zp2B�F�7����O�g�Sg�y��]�
�g�5�ߐ��Set|'���ĳ_c4ӭ��^F��{ ۉ�p�p�nQqY��Q�iK�:1+��􀈺Eȍ��y.w���yT�l��>tT5a�?��7��TKz��2G���5���&���HZ�GbH��}E���2�Ny3�'��oĠ)�K=RQ����/�s��s��WH6�3\;=�b�ca�1��|�d��_=�媮�ә��v	�6�N����)�l�5��.�J��/��y����L1�ݑw����������d��#X�|�*G�7o� �,31��Ř����[��f�-L걒/���i���</kF��`ԪWW�pS�} :�,X����7�O�c3����oPB��+o�/��#��	�B3@6_��yjo���#�U���i;� 2��EQ�?���Ĭ���T�6e禣�g-��/t�.��퍌^����B���Z�Ys%Wͩ��B�Tw|uܔ 4ŕ�S�W��׈�4,S=����k���w���/
E�E��6�Ay�y�m.O���yջd��gl]���R�(����f��ӭ\�*�j��
�:�����U�C �O���Uzi雦>L�c@�kk���K5��g���mQ�1�u�d�hCo�h�q�5_p����9K�S�:O���W�-L�=1�y61��?i�dQN�^}�]hv��Y�x�,G^/&_HP�)��k��ב��N	jN������kxY{Q��p!��Z�v����='�Yb !��@���do�{wG7\F������O��M��x�N�r�o8��(n�	1Lm��4 ���.�W3���/D����!e6T����tH�US�L�Ѡ��8�0���!�#�����uO���L2g���&����9�����Q6�3N�['V�S�Ke~��L���.�]yK ���H ��ň�~'��ȭ�O皗L���]��22fK]Q�|ǵ�{qE�xa���~N���ML ��o�\�ל����U�CK�Su�8G��x9cy(j��j����Wȕv�����3�i�F˃����Z[Hc�`��Ɏ&ɺ�^-{�5Ԡ���I�'�������l�d�f���o����-��%�Q�qK��ʳ%�ř#���@Z��e�#�γ�ޯT\ĩ�o��*����Ԕ��O%�g*�Y��تN2!`�B6��KٶgN�a:�W^8c#xJ9���N�C���K��C�-�\p+� ��?�5���ûJE��� ����o$��ؙ�<ړْ��o�I���I�B�,��3kA&��\�x���f(�~:R��¸���3�Tdb����o>	%\C�i�y^��w{ c�\|�� ɴ�?���,dxB��kN5Lic�����y�)5��<��N2���D����WK���7j�M�3ӯ�v������ᅗ[1,'	��ZS� q�M5	���S�������	�-ܼ&.ޓ4����}Ae�[�EJdJ9��ݻD#�-f�#&�V"N_u�1��α��F��M{Ζ	C96l�}K�o��Um�M)ě�vE��X"'���8qX�P���Gx��R�4��=?a��12�y��z�~T0c��C���7��>�{h�����C���VB�W����)m+*nR?o�}�hM&��F�!W82,�t۲����	�&5�˘*hrMň��^[��|f���ǶU��q�J�+]�m7���Մ8��I*(�4Z���*<3���G�r�A&8�Ӝo ���'>J�E����;�'�j'��7��R���_u����Ioꇇ���D ���]ݦ.�."�T�����E�T�5ǅ`��pm-H`P�a���H{��&�	���4t�H�aZ�K@� g�U v������t�/a�ِ�͘7����>���_"��?�P}��ҩe��E���iw�w��)쪧���5�R��^��_E�ȷ���Ao%�d :c '�~]f���@�z`gta>/�z���{��`�E�����($�:z��<��)A�e6b�=S�>j壁�y@�M~m��:�4�YR���n:D��������@�;}��c�3��c�����$�n%�����,j�I���3;Ǎ�ѵ�'{�F����I��΄�!MP�-�H���i��z�6ٞO���%`��o���٠	��#�`���o�0��2][�8W��c��O/B�_��.��7�w�3�
���x�N<$�A�e�w��&��� �K�h�;o�>_ĺ�����Ҙn�6�1h�?��L������Q����g1�n��+r�!Ni�2���#7�#���Mrs� �PvWh��&�ڂ�-3��l-A�B��e��7P��	rO4��b�	��RUi$i����yٸ�w"^������/��ӭ�"/���˚Q��y��~��*�n�7��qH�`"�I=�`r�,'9��F��Za�.GT0�E<H�	D����2�k	04�9��&�*�sǶ�B�����}���t��֤���%�\��>����h̺�'�<��''-�� �a�#qV6N9L8�*vZ/I�@�o��2��ríct�R��S����?8d禿+�EY��M� Z�gX�W'�&8u��w�ѰV�q�[�o[�Rv�>L�t�՛�l�xC�cǕef噌�itÛ��Vҽڂ֒�*�˗���1�:�t�'�`Ww����J���l ݍ`�u�h4��(^����$jx��s�~A�b���vEy?�=7p������ �Sݭ��B�D�ix+n���my� ����XW��<�"���q����������8���.�;��bw��%Uoɞ��vn�	��·����04��y�#��� \��|�a ��:���7���Ô��?Y�#��	o�$�����p�ELښ�!?|����&tA���T���t0�9t�E�]�mK��Nq����7���YFWa�� nC��lF{�!��<��I���?�I� �FC�|�9��|y8�=�V�����Zw�T�{P�x�R?�����xm�f%�Բ`pI��QZ�~�ZFE�����"�>��0��,/������q�i$���}CJ�,7�&���f��hp�m`S��tAPE�b��m"{pA���j��nY�
��0�e�ͧ{,�V��cg3��O���N�����<��C8�
�`������d�Jcu�Qᶶa�eٰ�9PI�*L�@Q�L�����a_� p�?���liƿ��]q���L2e�N#�����E>�0�˓͆P�2��5����~�4��V���&�*�֦��m*��입plʫP2��h
�t,�i�3:Ν*�r'
�U��#\�k��1|0T�NfG����[1K�ɇ�1P��`���n�H�rp&��FCBlC�m�b�3sx�H�/�?��k_���}o+@E&�e�X�[Ӈw@j��MSѫ��Ӫ!1+�����˻^��K�-w�3��A��I�T�/���w��{�"1��m?��;7�������^.[���E!��E��|��TX��R���Q=�{;���D��F>ѻ���8pÍ~f�m���}�(0%sfͶ�>g��U�����y�*��ȥ3:9t����X�G�Hߋ�i2) �Q�u��^�=_�*���q�Ժ�?M����*4�%��~^��/�wd]q2�~��l�M��f�[�mt�ճ5K+�#x@nթ�&��ǤSF~L�5x�J��K�\�et@d�-�>J�hG��ݑ�n�����i=J�Ք�[��N��4�_Jǚ�⛻�7	_�����w[<]!�&6��ԶłƢ��o���������ҍ���j=��<�RKIƮ���y_�yN8�N��	lAE�7�s�;k=榧��K	&��.�9`_�\4���7�D��s��R��+�~|���3O/��LQ��(�Y��>-޸[0�*�a�.ǥo�)��������6��(T���4��}9. ��S��%����#��P!�W��I���X���b-4pAF)��'��n(����%deRj�0b��
r$mU��9T�4�z�����AP~�	�-R���N�+O2���<PB���Akbϔ���ʿ���e����1����&��(뻎�@���NŞ	�{�o���(��_�ܰ��Lʨ�~g�W,�҇��	��ZvrE���#{����y�O���XN�<�A�^A������DJۋ4�R�:��<�1���v$���ఴ�Rg!B�ci9{"�Y���N6�/�d��;�T6�xBT|Zd�r��6q��]�f�xf���%Fʸ\�ǌ���`�Y�ko�����j?�$,&Uҽ��Q�|G:���OlJ��u�B���Oe+���k��)6/6E&�����Zs�--��gD����1�;��}mY��gU�9�o*�Ў�J|��)�W������qG@=�6U ���2k��w�'�bY�Tp�nm���p�X	 3���m�,x�Q5ce��}o�l�k��x�2PW�A���XP����쯴���tIn9�@�p��3.b��Y�Og<�S% �ڦ�C� o�N�ͯ�0R�}[k�s�l>�f}�q5'��s���*��a��T'�v^�u��]P�Ö��z��N�f`���P�Xw�=��Ň;a�y0��vS���T���+���b��D�>bC��O�	�8���bC�Ȩ�d���a��zs�2w�wA(��vXg5��<�T�*,���,���5����'�Hh���L-�=��� H�!�'�_��r��6�RZ� Z���8������V���AzI00��{ਲ਼��o��J��_����Q�#ԥWX���e2�g��[�5�GC�^���#x!���/n.w}
M >�>�?�FRR�&ua'��{bk奄Y!s�B�h]F��4q��ȋ�I��:aA!�*��d��3@��j@�a��&K�م�(:z���։vC���|������a켈a7�|1m��y1
TI���;p.G#���>/�* �V�~k�����g� K��o��ƍ�Y�QX�w��[_F{4�~�>@IU8j��蟤�VH| /����|��T�a����1��cS-��m���)� w�!�G����f�Ω?����٧�b�Um��sG����ii� d��C�r����8�Z���t��h�p\�G뿍j�=Ӧ�eT$J�������?Qc����gk}/}J��6n���2%�步����mǔ	�cc�4���}Â�}��W�3���%Jy�������#~��>N�;�N�2N��������1��M���3�p��ߝ�[�\(.���|�X�/��Z6�K2�E�J�JN/�Y����E=�d�(�"fe��5� �����s[بm��u�W��q�i�Q��w?�Zt�K��]^'Ҳ-4�RӼ�>`�/�DY�'m-T"���mT~H{�Ȯ{�&wo����l�g�2�=%�v焉vb���N���ö�;��A�KO we�%�u�"{�� 9z�E���B�����25�}EoޤO�@q7�O�>�z���h���R%x�,)O�L0����
Ŗ�^�m�:�_�o�>������&|���X��B�=�C��L��^������^I�c��Q����)�C[��kvn�C�����ȑ��[���J>%����c!љ.��&2�K k��d4���n��Ƚ��U��-畑\!v�0��DJLk�9$�֙撪���O��.c��.e$�,�rm4��B����`�A2��/�����
i ak[�g�7,���,�xy�=�#�r�r�'���z���T�,��s�G $hƵl�,{Z��la���ɘIl`vG�s�Iɭ�#������*67u/�C�!NjxV�Vp�v�-�&笠��ls|��)� a�I�4M,'��[���g���Ht�d� ����^OaI: t���y����a({��Fɯ:>��l75���N�j�5���.B�h�ė�*�f�|Z�)(��Ţ�`���DoC�y�����8aIW%��� Ga����cWB��|�ix舶��o��G�9>aa"�s(��L�J��LU�qP� -G$��ku˱�b�	�w�[2@T�엧��5�tW�mg��K�EGq� �Ӆ��L����;�C��U�-9":����G*'��S���fk[���:�"��V@�e��(&I��L�=��F��FCl8<�TK�'�����q֊����!�i�V�O2y���R�~� ��V�д�X������6�� ز����IHlK��Dʮ[�����2��-8��A�)a�Dݘ���'U1�[�{ݍ�Ջ�ݠ�m��ڢ������P:y;]m���]r���Ny4����x�T�E�b�1�m\�{["E>�;<~�V�\Jn��_����`��+=���`z
�mN�a�+h"Rˠ\~-�/�Ȓ��H�?��74�B��^t�~vB��0)�6n�J�	ml���?xγ���D��XRA�����b��eo�׃�6�~�I�����' ;�}kH����TT�+KH/[�s3GxFi3��|���������J���	����1��P���%Q�3�)�=�7�E���.Nl9��������հ/�f�Xy�I��KˀU|C�E>�sٿP�c<,o;���=�iY��^M�b���i�zgB\����~K��F��RVU[f����)0^QƶϮ����/�bU��������Rd���M�WUn�.c�?T��L����2�3��� �
4��@E?]��������Ȓ=B�~Y���ɺȫS�����t���z������M�,"72W
��o ���$�E|lb�h��+H9�@;h*{ʫ��G���kԱR@���]��6�AKzN��Ec_�� �3�k�eo���`���sC��E����o�S��w�	���ؾ����>s}�'EC�aAZ�ʍ"LNP:��1}?N4��t�2�0��x�"VU�/a����4�t����ً棼��="D���H.F�Q*<�˿[n�w���8�լs�D�]���;kp��O`��Ja;z�7Ӕ�N4)� c��U�����g-�ڳL���HU{|�Jc����a֋[�rX�f��~�1��k'��z�QK!�9H����n�(���.�VQ"Pf�iz�ZZ���������^����Z%��C"r�Y���%�%*�潩�W����L��7#�]�ݓ[�ś�=e;�v��������2�(��@���e�	.s�
�k�Iư4!�)��`ӟ�t�0��*�C#3��]Tn(�v˼�z��{먐|F%��!'e��}y���V5L������ wz{�t`3�Y	���ܐF�A��`�A|2.^q��hӿ��I&ep�8����|�K���,��( C�����7ǥ��bB|ڮ_�h�
�s��uI���l����ᾳ�4�P��= %_�HQu+3�1��C�P��T,6��K+rs3C)���u�� '��CN(Ĝ��2(�6W��q#G�M�/�n��|�ނ�v�d���Ċ�I�b8�y���G񆚞h'�H2��ׁ�`��yI9��Z
K��>��3n�&A��s,�?���gGm/lEKC�#�5#%*��Iؔ�;��K�W`�3�~��+qs;��F�Ô�h4ޜ �ej<b�̀�����9�Lլ����#ID��T$v�HR�K�712<%�r�~pB���X���9�` V�@W4/,*]��zT<�7�~��26��!<�z*2q�d :D����_����ڃ]��6 QԤ��ܖSs_%v!���k{�W]R%S9��Y0%��Q4�nu����A���v�A�w�����A}q�B���`ogO
CwrN]�hZFG�O�o�}C���
2��r�hѼw���[%�υ���3u@���V�Po�V��N/�������nm%&񨹈��VQ*��i�JB(��y��� ������*�j�u��<��Z�ޙ��Q*���XH��wܯ�_�!�.(�G�DOwX�sU�[�[ Z�Rغϵ�3-�Bf`�
����J��J��� ���<��U��7�
/V���ۀʚ��*��-eᘡ��y��ͩ:aћ�;+-�A�Ʋ��.5����|���R��G�Z��M񴸦����r'+�<z��t�V�8�L�и�~�f����x����
�D��*�9~9�>,_󶚷$��{�>���9�M�#	-ŏW�\��?�V:$�p`Ϧ��^R���E\�g�k�$/�t4��W�/8bڭ�����͆`^�B���U���${0�����!UEd^e����_kb�F���B��l�w�슫��I*΄��	Ӿ%I~�l���� "����ia���DE���x�����E�b�4�8�w���O˷>�H���'/���|n���[)̖���{�7�\fy>�S���|�ޞ8�3�_Z���܅Os[��w��K .����]UE�����>A���i�[�l�&���Vm):3P����]ț��k:��,�6����(H�wj{�-��QH6p���d1�7�LD��=��}f��JȐ���G��WTa]�^w�G"Z�u���������3����Ui��*�/HY�����f�ˮ�`6:$c���K7`/`���Z@9jރ�Ũ�3�������t>�R�⁣)����{�>o�Q��r�-��>�WR�t�����]!�^�[�sa�۾d�f���}�f#��(�y}Is9KG���;��+I{gآVE���c�ci#�YkI��{���l��굗eK�5V=>�'ö́�os�XN/�
�k
}T�n�Vp�Ҽ�%��@t<>�cdLy�WF�[�$��ij��,[4G��/��G��/R�3�}�XxС=`�cO	��Yq�}�'Qs����G��7#֠[ݝ.B�p�?1�n�e�a���q)0��������m��U�=�7���?F�����m���_f�g �J�"��)3;m���'��M����M&��&��21x��EVt��#=��?|5���8
�ːk��=�o���ɦ�fx�B5fxV����ș��B3���{�=�E���+�N�;��l��\�m����j�׽��!��=bz&����8Z�?�G�w?�����|��:?�r/������G�U�=";��Ɲ���I3����7��Y9�)y�;fv`�%gà�e�����]�W��6�
�D� t�C��[�` �+b�GW&��Zz�"w����e���M	?#)��+��b��m���N[�N0��`���oG��1!|8��S�<D����#)��w�����������g#}d��-**E����Ɛ[��2�d��%f�V�W�G�%�x�.���}�u��+�� �g��G�ڏ� ��8��c��LF����ُ��'r%wGp��Q��xW����4Z<��h=a��E�S��, ����3I%����x������X~huy�϶ ؄Ļ��c̏=�,���W�;J����6F�e\�%����^�9�'O��p���녔��5,��N��+�R�P�m�Y�3��ҪϬ�3ۚ��3�����m��5#�w��xC�����}��74��/��m�~��L�h� �U� ��V%;�#�a0F��wO���ؐ^�72{)��V�t���h� �UOȟ
��V:�#�*��N�-����(�j�.>�h7K`�O4�hL�uV*F�$�RA�����;�z�RH��
0�$9�wdp��oѰJTNE��G�R*d��(��( �ݫN��MV2���9og�/3��~.��rƼ�yÏ�C��FA��:&�w�(�
�K�+3��'6�E4`��R��V�W{Xr�-���36�oT���=��j�	�VױcQ�,B�}���W4)\I��IZ�0��=m���}�<�	E
l��Z��8��%�ʑ&�Ȯ&8�c*Z����)�9��Df$Ҫ�Ih��S���뎨���l�7�`m@|lF�y�ǭ�_F��= �dq���>�_Ti}���b�H"f���}�Z��1���`��y��h^hK�`�zR�$�cʵɵ��@���%��H�߻b���gW/|<^<�g*ʬ�(�^�e�sy[����� /g>���D.~���p+l��(A;kpT,�D�#��h��T�kn����C�{i����ai��~>[L~O��/x�1 �,Mj�̨y�m.W�Eߤ9ԙ���Ĉ�p�5�Xm�H*������%p�M��z�0X�$�w�!a���A���W/�vD`3^�<����i�"�D]6S9�7Jn֘J�W$d�T͑y*�4K�|
���A>�;�"Ζ*8����x��Wk���Q��ǘ4�s[��R�;��x=OX:��B=[��+�g���LU��a��$D�5��;��!y��u�D� �a�:ćӍ%[;��S
���+���=c�����6�a �&� ���C������"�q^����8<o9���M�0~@�л��U��Ƿl��j+��T&�B�3�
�a�#�~.�C��Թ�����jF� x�e��#3ۀ��{
��h].�3�v����Z�5�X>I��0D�6��JeP�#O�xϥ�޶��:���ɼ���� 4ģ1�	g�ge�ߡ�#~0[-C~�J�69:��B��Muj�U����"�9�uowS��;�~3��绛ve���P�M�U<bb�*��2��YQ1�k�G�u��T\GyA9:�I(�#����붋/�}�*�uF�n���i:ĴѶ��o��1H�5�5f/F�}�ypT�G����Z��/��
�g�dm=J)�UG��D���vv,�*� < �������0���<�b�-��>{�<��vS� I0�2 ݐ���,�i�%��c���~��Wj�8�ϣ��U�p����GQb��;�����#^�5aUW�HV��{$�6�v'�"��t�n-�e��3%q&�]ݕ��,�V�mL�򮌋	Λ*ua?���:��@n�q@������k��E&3	����Z�^�)>� ��Ce'r�����	�w1K�1?T����;��M-��~���T]ky@�3�$�L`Y���MnXBx-b@K������	\@���@~j�|��m5>'�
2�,88�����j7�����W"�W&$��2QsQZ{���璥�wh K@���)���%Ŭ4!�~*8�h�����%�H��z!z����t&v�������rg	��/Q3��ΠH2룃m�	���De�Ey���H5��,��Y�CŢ�����᳅��Q�`'���6z�K9F����=�)����x���vR!�ZU�����"`�/h&|��0�3uJp��&�Rj�,�U��j<���j�0�.�	 H����zM�H��2`���|x����)h���Sh�VQ@_�#҇(��ePl���"g3<JW��X�i�����
����%��p��ᆶ����Kh0�쳵����%�6��s��&X�Ep9I��ޜ��H�-�G�zu')��o�~w�0�] Y2L�֘!i�ָ�>J��Lê��k��d�f��W�oRo]t'�����j�t�?��x$��ل��p7n���]��"'�:��������=]�Jǧx������2T����*'���
��W����燻��W�U�yZ�!%*����`ɗ�th.��B�j��}�Te"N�B�Hs�ݛ�Y��)ߣ�7�r ��L�PB��m?�d;�V�����Z>5�s8᷍�~��;�_�e��r�qi�e����b :-�V���]���:N�l��5ח���a	M�X �@31V��,0L�RA��yxwm�_�B���y\隃`��� Q�w�~QW��'#�#����0|�w���e�z��QI��}����fp�x����*��+��%�ݩ�9�� Bӎg��E��j�梏U�����^(�U��$�)��V��w�wjPƙ~�b��;��*�
X���5�f�^�;�=���E��A�8��P�S�QIK��{0�_��̋7H��R���8���K>`{#:;���E��cC��F��G2�ϦhelM�@�Po�U�oSEY��ͪ�g0;/���o�7���?����^��F �A��:5@���q��Ȏ�g�!Ct�hL���nF|=e{�`B���b!y�Ȑ�<�QV�2�q��Ŗδ�K�����Д6�\�����<�H ��-����W�v /�2�C���
�x��7�Q�� �x�V����gc�X���M��޽'�9���ܧ��9W6)=*h¹����qx��Ӷ��cUu)R� (��N�nk�K�c*���Xv�hb�G�-��ʦznA�ă�a�O��)RM�6X 
d0��tިA�T���NH<QN�Z� ���~��FU\f-�]�v B��Q��,��O3R��6�x'r	�8&g~C���.��ی׀�n�&LR)8UsA������%�a���)�lb�+�mfI�iGP�&���j#o��1O��oCh����V<,2�|� �IcCK���e��_�l��t���O�����t'+'��я���g��m~�t�4�-�"<��ҋ�[�9�O��O��"M�u㠪��ڀ��ZwPr���� ���s�I\QZR,�ғ��9�A��q��5�g �'� =�t�H[��*Qp���\;�ȟ���,�É��Fڡ��Nf�S�BU 7���PWLs���(���p�Y����w�.�־�]�rY�����2J���6]F��-�^g��7W�4e���������t��(��Zoz���FC%,D���B*n�Z��Kȹ�/�ԡ����aH�Ք�◍[�=U{��CD��P�fR����m�>Q/��?�Ir����N��m¦��Y= &-��BQ��rC:����k]+y�]��&�d��F�+ߔ6L�~����S�"�+a��4k�6�p-���]gv���2^��+5O�N� ��;3Is��B6��$��8�'�ɵ]�x�jO�3�0o��=�?Xd��.C�:�d��	� ��L����_���B�M��Ml��M�)@
�����X��4?`����y���+�R��� ���ݍ ����t!����;ј�:��C�B�g�*�g�W4%�혹փ�9��%�k�4���X��0�6d�W��rH�`U���E��jV�����;'h��/M��||�����P7���`=U㲚�h��XO��s���$�9'���7E�=Us�zXq��5�pi�DY6�ė|d|����SlEGq{����z���Pg��`7��as��^J'B��-g �2g�/�;T��
V5�h�hT�:u��Ro����~��`��0l�[}%'8Q-�����P�@�O1����u�L�'��:Q5�W��YR����ف����o��D��p�����Ͽd��6̐��d����w��3㤛�n V,N�:FO�U�i-�Ks���6�<����ФW��Z��e;u�sI�Ӳ���
[b�30ͬ?V��,��=��uz%��*��t�5���lP�WHΗ@J�̞+|�7���^��HO
����uO�o����H>+X����ܟ�lƉJs�A4ocΥ��?B,Ӝ�M(�\��F��A0��D\�1�P��oE�M����%u��/M���){F%i��?�ޞ�9�C���CR�z��s��&.Hږ|�NV+
~���~���������"Lf�
�u�WWEd�akխE���r��a�^��
+�c��8�6��'!� �����p��RąÞN�V�|r:�#����V��!Hl��������=j���'�6EY#��C�P�-(T��0�m�����@�Ӿ�X��#��7_�O�$Ȉn'�(YP����Q��NC�*v��ݣ�wT8V7��:����k�R �ś�d����

7y�;�U�T�YuEh�-Y=n��L��N��-�*�K E) EWpM��xv��s��UP 	G5D��v�-�	BY��{w�N��U}mq7	/㉄NO��������b��f���$�n�Y)���
�s=���RV ���~!M�?���{����c�7:�[@��|ؤ`i��g@��@�u�}�@�|}�:<�hW��V�z�gֻ<�d��<����`Z8� �;�W�	�">lz�3X+ʚh����i/p�BP!�d���M�,��,�T�3�&�`&h���O��ñ��v��a�D��P%��ѐ�y�K�-Pؔ�i�|��e*��;�X' V�F�dKs3�́��tM?x�Հ�BB��ļ�u�G����q���T���afx��.%�g.L�J���#�?'suƞ2���ܪ ��Y�J��K��HY+c8aD�V��F�?"y(qq\��H9�T�S����Z3���ӱ_�i7XG.��j���c^r]����i$�r{z���Q�W)f馈Y���D�c��Ĝ�.���އ����!�	���l��LgǇ�Z ���Y������Wd����S!}₁2i
<��=��a7�C�,U@�`������Y�L�b��c݅�]I�ykr;�-H�a�<K��2[��K$�i�q刟@�^12��z���7��9xL�Otq	�\F��b���+=Nm�e�D�^�f'��*�{&c�"�Hc�K���A�
LI�ɚ���Rw�J>M+=� �3d��ƷVM3|��/`aH	lE���e��L¿j���)H�G("�ë��fV_�:��C�h�f`���i
u��C_����2�Ipt*�>ڐL�#�������,6�M ���FO>����x+�"����U��,*n�Ի|,��f$4�H�c�ҟ��
Ai��Ux����V�B{�B�7M�8���)#SZ���Ic����:i��C��J	=�o9��bj���'�؛ ��t7��*�����FH�J�J�r!"�*�sV�X��tT4�2�䮨깅
���a[;���L$I0cD�Hj|�v��d�4{eP�˩m�ժ���{D���/�ҿ�����J$5D���+����.АBVP�����H��0p`ތ���@~�ϊoKsΡ��0��S<�<�sԛ�SPF�&���6P�"j_X!	��O�<�+����ܟ-��d��Ҽ�/S.���>5(�"�?�]�']��K�U�"v֣4�� F���VPkע~H�I��tq#_�+� 4���-��݋�p�dA����2��h��bu���S9�����jZb]�B�A��QI:�j�$'�=���j��f���U���&[�U�F�S�5��{�_˒��g��7�@��I�`}���m�v���W]���P������Uӈ�h�����|�
WX�[�opm,!�s9��'�E�]�S��r�wb���-�����q� ���,�cŎ�|g���D�w1e�+*�̷�Uw	owA0)�l4�\QRI@�ŉ�%��[�l�F5Y\�4N�§������ t�w�ٟ=���RK6��W���_\t�����g�0<��n��,���flO�I���dpa۱S��K&F\k�鸾D��"���S�T+�k���� X��M&�cF0�$x��C6*l�=ݶ-��n�A�h�5Թ���w�gϊ���`9��Lv��'o/�ܖ�J��C�f,���_\��zA�a\�m��X���c%JV���J�]�vWm�6�k�c�v��L��$����i�e�5n��;j���(c���⾅~�go�*����IH��ޛ V����얘�� ��w׈}�}�1,H�Xg��R7��&�8��Q��A�W���Sc�-�{�wXR4"s��6*���^��9�*�3k��L@�NvҾuT4`L$B�,��rgEq�m�>���_���w%�[�T����!誮"PY�$*@�L"�t�e��)�K^����`�\��ۢ}�ֲ�������(t�$�o�^��uI�D�X�5\tXW��@N�@�bh��B��#���?�n�k�&�Ō��2�)�~5�D��{�?���РZ�+$3�j6��g������JW�&�ڕha�GU��D~���T�c�ˊ	l
}��H I�������L���@z)���HM�8�e�ҏ�*\L�o�
�P�G�֡�k��.ҍOƏ ��f�i��M�F�j]�ǃ��;ܻ�R����x�6Y�F�Te�eq���:SЌ���n�3���W< �UZ]�:�x���^.b_��T�}*F�R����1�鄈D�����٬�e� �$���b��7�-j��l�#,{���L�s�hQ��tɟ�Q��~�[��+ט����|\L7�6f�[j�8u�l��y��ڽ;H��'β���ܜ�� �cD3��>i��~��t�ʱ�2�Y�Lк��u
�؏����H��ٌ�P��s8 ��[R��k��z�s�H&F�����ZsK��q��S#��r�
�N���t�nh0�2�{�.�pܸ��?�a��p(����؛�˛�'B�H��\��p!Y��Jvp1���s��}84dyv>݇�uK���&�����>��.dKX<C�����듸�5�3����
L�穰���ӱ$�C0��3����9��$�]~��z*�Tj��'�n���<�-O�����7^sW
��oi�~ƭ�%��)%	�qQ��|�8���O�淃lD�g���t�ii4�=��-�m�?5�h��g%�h��a���2��Sm�A�)�N���w�C���K����O}~H���-�6z����OR�I�ߊ�vŨt����%#>���U��8>N�5��V�/�>B?I��`'6���n���,�k7���y�]�P����2q!+��Θ�V���-�q�M�Y���O�m�~��˭���2f�����g�F w�g�f~>Y=�4ɝ�+S��>���X��H�����{4�+ʎvz�Y�D���V���u]�g��i���~3���_���l��rG{f5�95f��*�OY��Ѡ������

9�误��{ҏ_LВ�ĨE����>��inv������޶k[�J��fW�������r�bv���"����c�
���@T����8G�w�,n�k���$���T�{CN���Y��(HZ0̮R�rn9�{�X ��xD��s���*�p��G��p@���&��=�m���M2"(q^w*����4�i��(�_�^�У�[�2A���c��߽x�uJ���ۚlQ���_5L,T)�����o]s��¦�|���K��:����啾�\�k8��џ(
�\�10�QL�����k/<�C�ѯ[O�W?}|㧱�|t�����]�A������w��[n�$�`߿�R���F�Ս|��_[��l2J��!,���d���f��o&[o�e�����|�dNG� �Y/���:��e����k�kJ��X6�\�gF���r(��toP���	�kZC��Ӽ�FN!�h��3evZ
>W���6�_����6��'o}X��sH�8#��_��G��$��7�`���?�pV�m���B}�(�y.M�䧓Q��M6<\��{��ˆ��x�Y8If�g�qO����o �IF�H��:;*,�=�1��j%�k�a�����������
xϴjqfه[;k�9<N�^��s���	��k�F��J,G����½g��k���T,����2��Z?!1���/���
B��doȯL�h� UbX7���"L�pPCַ���G����ik	�|���4�VX	���z�l�4|�}mf���ʕ���C�܂יּ�ۍ��2�-J��C��cA6RXg/=�Evw�T�5�����r����������hŽpgqyl�E�=�{}@�}�8I=��`��l�̘�jz
�����.��,%an����I�s����L�ϓD�g���[h3�yX�+τ�4�w��'�kw�"$Q	M��Xi��m2�Y?�l&K�l�p˳��39�N~���,�E�Z�t-d��
̙#��rG.q-[�a��&(�Er�g����{J���L6\,�c�q�K��i�|�MUBR��yy��&���mQ�b��Ksj�6�4	��YH�KS��:��v{��O�>�i�o� �։5�d�ʍ�/qÞ"3����-��I��h3�j�r�m�S:�YO��y-��؜�8K׭wd`�*�?�q����Z�ZW�W��xU�b�8f���[�d��뻾/��͵�����^{�-����ͼ��H��~"E
()���@�r����
���>�z�Ԍ��oV��P��V��?_��g�������;��JuI0�y��.c��kU� 4���Y�F���>���/�c����rFw$��s��S���Y��h��*���҉G�4-�a(Z(%l����Ǎ\D��|M}<f�.��o��;�͑�8Ĭ�͜�<2��
?�v����a$I�nȯ*fF�����71�rM���Ǔ,D��u����r������jc���;)
v��T�l��(ĺqs"Y��b[لѩ�Ҵ�N�m9\����}v��A#)fA$��M���Ot��R����5S�+�V�6�ɘCV�#��X��h���{�R�%���s�Qn�sXI�M��M#p�-t+̬��J8 nzvLƵ�=I���4Dv��"xiΙ}�i)��$�
C��J��<L�u&)�T�0M��l!�<*��gL��̷{h#M��44��'@y�a�.r��X/OZ�9����6sY1}uK��\Q�)Z��v���2:�ƅ�.����Y� ccW���7I�V�+�)��?�vŴ���cB,���[��0Fw5�/>yi���m|�s�kI�FP�ʩ�J'�r��*��r ��us�K[��J��=��#�Sx��q"�6;e@�ʀ�{Z�_��;@*���N�/���PhT�X�,hfK��ܗ��C�I��yСq�Y�l�G濼�_s���c��P'��g#��>���Y�B�'�
8��w�r��Χ�Ϸ���v4n��VL�7*�<jG����Jp�Ɩ{��*I]���)b����z*_5yF�[�ҭ`�h�WIЄ�5�a��=�AI�'3h�vG���B�?�_�F��I���^�|V�W�r.��x��|w�ʫ��0���d�'J��([q�XT��(�ҥ���O�a�!���w*n
=j�o��{�ҿ.��ɧ�2Oہͼ;��\��6�������)�4�+շ�k_�:�sB�L����Y�2^G�7G_];�*Q�;j����뫖\��o_�'�����t9�c��2��OՖ.��k�׉�'I���D�Z%�l0���]�W��3}s	�"�([E.@w�`)Gs�CIc.m�5���Ѿ�����Gr��j�P��%j��r?��8.�~�O��Ǖs�$��(��-"e���\����h��67[ܭ��q>��7|�k�{���̨L��J�M0[*�ճG��^h����C����l��<ٲH�s��KV@/��Q��­T.A�x�H����
\m�%���k��+��n/����<gZ����~_�S���-��
�&���q��N��4�g-�^��`�j��'Nn�.�C<�C�Л��Vh��i|�V�h����f<�ۗ�n42�j�},<	�"���Zyp�t�Y���Z?s|��hyY���*��d� �j9@Mf�Y�yf%U�e0�$�~�_s�?�a�?$��DہY��Cgw��-ݟ�1N�����܃�,��T�������D��!�G�]���IQ���O�.5�i���-	��&���F��H-��l�F�@:p��g^���{5�d���?[l��>�X,t?�J�r}x���=��rل�����
�	 AC��3�sl!�ؕ���Z�R?�_�?^�#lgYe~�I³��xEq��n$Q��d �C]or�g�<N�\)9���\��d�ӄ.v=`�U�����t��)C������X�J�
�H��
��A��e�A�E��Ld��ӈ���>�" G4�A��r��
 j�~ǝ�E�;8_��L!H��q��9�q�é�-i��p���FX�~N�?A����WjÕ�8t~2^�'�ZB��S=!HEEo�g(=T�X�k�0�!<)�"��N��AM��0ܭ/�g�{2�%�Z��L��NZ���]k��9�'5LC�o����|W|-?:X��<o���s`�#;w� 7Zz"�AL^�䩅�	�'k9�$x���Y3�,����m���6�4s�&�AA��oy�!����5AJ}I�ވ�&��]��|�щ�& g�-�my��A�c"�����D��0��))PF�Hڻ�Zr��4����ʮ��8k�Q9�B�
���Q8����AT�@�:c�"i/�2FFy�9�A���˓UQ�R��Nݗ�odV��N+6��ܭ�_G&/����2�<8�'�$�L<n���k����94��;��7�CqxC`3Nb��(��ː�*�ā��x����5%,ёđ����Y.<p�<���z��2���e�h�[�S�/!���"!i%K�J�m�?A��^ ��X�-d�'�35I~� �t~n����T���c_?]t��w�4����Z��������S�lcL{��)uF��)������їQ�NVnx�9hB�������N�#����) i $,�h/�M�)��6���	3����T5�)���@"z�vO�~�x�Ou���[4u��@��_�����k^�;�My*�8a�	x�d�f���ld鷓ś��>??���E�L�_�K[�F��ńLC�s���>�-����Jc�fZ��1�Slo�B	1xٺ��r�תy,9AZ��HS���'����&V���w�~#q�lx����=��8�^m(��A�s�Ȅ�G@qjߌJ�+G��w�]7�aⒻ3��8��q�($򻊤�:^�3����4��|�N��ڞ*���ЌFr��S�Z��cF϶e�C��
��$�v��:���n'�P)L�b���b��7~�5֪\�ͱ��r��s�n�߉�V�Κ��>o� �ÒX�<�F�&:VD4e�=�?���� �ƴ�03h����\*��u.�P�oB�I�Z���u��t��=������"��ᏽHE�Φ)^������;���F0��4���ld����Ӟ��{G���Lˑ<نh���mu�]�0��
Φ�N���1޿��á��Ï�  /�ڋiz���a�%_�̉�%��sL���k��tL��X����T�?�k�钢hqV����O�r�e�N���+K@H.�!�>�g0o�پ����.���2=]�:�]���2���E\{�L s�dh��5|n��An��m_\� D�����w+Hz��*��`����s��b C� #
�<��a�dA��us4 ��_��M}'M�륷�t��UA>�H��B�\�TN�mxC��|�3}��\�`l&Ƚ~�j��II{��^��K��N���{s�B<��������3$��hg�EYK4E.��h������l�h�=I"
}q�jʠ#�=���=bA��"Cƻ^��,�m#
��Z���f��Hޠ�H�-Y��F!zk�"\i号{�4:�
���礽��͜DQ���A�>(1!06j1�&����!�e�RY�w�Y���>���XX�wk׼ ���$�ٷ6{W+�8��<�NKQ�i�`!��ˇk-5G��9%M���쒃�瀹tS��-0��J$g�;�uv�s�&�,�����ĸ�Ȅ�.މ�	��$�[���՘QD9���俰i*I���b���2.t�I������ۡ�ˀO����`uƚ��\)/7'�i��_�8��͚ҋ�$?��K@�I��GF���>y���Q����F�ty���ʶ������{c�ǒq͌���f��D���[����
5&���i�.�=ˀZ\�*u��z�� ���=%�E��X@A�L+�*�M��K�E����P�c�@�M�(9�� �ej�%zq��a����8
G��!�����!�V#���Ţ��F�r_]�o�������S�-{�1��,C�Y�#Hs\w�LG��`Q��w,\��q���J�j�p�;0��_��<���p�ɶ�T5V��� ��4	�{�r�k�/�K�������T� |5����!Gr�w��	OMa��&�?<�k�@�*"y�X3!ށڵ�GZE�o��}/H�]
IT��92"�����ؼc����r�E��O֞-3�
3��m��������aƭ�����
~+��-�y[á�b���J$�����(��e�(�4s0�mn��Lg�c3���x�:��ԑ���3�ޕ�BK28�N�U�m(L4�~/��<���h�̂ai�|������K�����ZQG�,rj��s��У=�=�<>A���kDc)о[Gۙ�1���G�=�)%a%�2o���������bW�9��B�)5�\�Tz��k�Y2�Ϸ�� ;���g���M5kzKowb�����`QFԫ�(���P݇�����O6j6%��>�u���z�>�Sou���>��쁬�L�`�����O��ڼ�u,��4���Q]��g�����/ܧ΍,��?���;�3I��_�Ѯ�E�*�ւ��T';�4���Q�Mb4��&#F����*�l��s=3�T�>&_Yv�LQ%৐HZ��laՐJ�8+VF�!奈�q#�TH@�u���Д���"�	������'�� P�d
Z��;΃���B}�W�D˫��oK�̬zb��˲:\��XXL�ƂF�?ՁcLU�^�50!*Wn;��6S�`�ܠ�#=�AŲ%ck����Y�O��w(��cB'@^������8�p��lz�ډ��V���Z��8���,�JyapY?�(��`����� ;8 �0�_���
�1\@M�������~�4�W�0�8���?!�rHX� ��g��' �?=�(^�����d�0��lg�
���%��4;�R��˓+
\���{�q� ����2�iy/�X�6�;���bD古"���/�t�G�}�z���*��/�9�#p�]��w�oM� 1�J��}��`�RbRzul���ڋ����r�ˮ�z	���e#�}�$%ač8�,�p�VӢfU��S%��G�Ƭ�`!�,��m��}51�� ��<��P�a��,���%� u��ZDS�_�A�Ӝe� _�b��A��L�k�NeW�C��������Z��f��j�B�Z%�)�X���j6���kyc$��w�߇�I)N֔�^�I%�h�曱nf�tC�ƾ��[?�ⶊ'�+�(�Ӧ2��!�h|��;\��@�$ɮ�V��Y�:}�p $�;�$A��N�q,,N�&k=:�r�gK���K�f�H������
� P=wj3��ћ@y�goA2�{��E� hH!OVe/-�G�.o�q��#�'���ve��T3:��ޤ�yȵ���O��b��^�Ε�F$Tz>��0i�����������޿~����+6gq�����
�4o��|���׾��y��pz�E��%���LS[�d��lH}��{+�q��uͰ����cS��m�p��l��%���f�| ?g%J�X����ׇ��@��:��7������Ͷɴ^p
����rD�����������
�_V`��~�����.w��v�Z�'?�j�;K�{��ka3���/�b6��3�>>K\p��j ��?��AS��7|�RZ��(D]n�/`}�CN&��]�\��@�6m�����{��<x�D�e����a+��[͛�����>�J���Z�&z�Y�-��_2�UG�'�yX�������}�ϸ�>�)��@�=�(�����v9�iɺ\�s��:�~n�ȧ֋Ð�g-hp���^ډR���OI��I_�Ȫ��"Ig}�S`�x�^������_6p,ݥ:�d�֎�_~F*0�4,��|��m�n\o������MyՁ��N��Yv~%S䅍?壔)���ܤ<P�m�f�-F��K�/���	����ޫIDh��0��h��B*�a�Q�op����R�L�G1��d��G�--�nX��[����,�aG����Ө̀"VP�\pw���bꌟ�>�fK[Ɛ�0įd`__�fh�C�w�q�I-�Z�z"�ȱ�þ3��<O����-0Slg�gJJ���8a"��v=)�Y��E���y ��Ǩ�O��a�s}��D�)�WY�mz μ1[S�z0q�����-��-e�:���FG����O��Ι����)��S�q�f������Ɛ'IK����O�w��uJ�/�&���4-�6s�⧃\L�g����oƼ����\q�5ޞ;�i����m ������/8q^�us&\�1�֝<i�լ��m�m+X4�?��I��R��Z^Iۦ�녖��A�����J���#��������빸A�Z�ERq���"r�C��,��0���j=�c�ȣ���O��3���}�_���O�T�{���BJ��$5��
,݀I.��M�vAn���B~�2����.��n(EZ�O;��mx���t��( &K�7i��L�`yl��f:���; �n�vE���M���9��>��C.������0�����s���#�']��<�,��b̢�q���1���y�e�1S���_=�V��ál�j���i=��)�ە��?���A�px��uK��v�&���Mz��i7��x�ġ@�4]��_�E�K�3���8�]�tVc�>��'VlN�Qd���k�?��)������J�&/����91�cDdכ��B�����*�k��sN�a�۾�+Q�rc��aӲo��dYpdw�i�$��,���
���+dSj�kR� ����F��Z��x�2t��[ʒ��$�<2���
r[��#���9�ǽ@���em)�ד�����,��u�(����W�&�_<1���c���:I���Yt�ʘT�a���жR���6>�Ot��jpV3cخ�]���j�Y*�>p6vN$�w��V�b����{�6�@�l�"�#�[���I��*��
Ď
��O�V���Ou�������:H�3�ywc�=�[Nh��O_SR4=�<��;*���N��.��P�.��"�C�1�Sr|1�R�z��h����{�z���p��9E�o��jc_���q�)!�lr5�w��#E����^f��|������_���(��֨g����;j�rr��@ Q�M�}��J�[���8i�ia%F�FA�	G�}r]��sQ��]:�h�5l�G��H�K�a��|�Fj�����$#l�Ae�˷�@��:%p+�yϖ��j'X{<P2X;�tݝ�e!P� c��R�.x����wW�Ͷ!Ԯ�W%;j`6��s`�T�`��� ����	Y�g4*����/�ֶ�9zŴ��k�=F�Ii��`&la��k�̔�Tk��X}�l>mAzw�sW���I3vl������9��Z"c�J�w��1�G�?��c�m�����I�����=� �U[�6+�6�QQ`�	Fs��A��E�6�aD��?�p{�oخ�2z��s�E���Ȝ������W���d���G�W���}��V��\�1�̗�����~݂�q�N�;Z�4�ǰ��!X�6����6��j&I�ŵ?s8>1Ңo2�[���c��Roʹ\T0����6���r�6�3JL�P���G�ʫ���vӺ���E6:�4�o��Lm�Yhb�pal��˻��d���ێ�,i����S���78�r-��Ϻ+�Х��=��ZIs����:H���}y��5C RV��dI��ڿ�ش��w��9�����E��~�-@M��+�U��y8���#��o����� �M+�f��M��~�v�1UCּV�mmf��T�Q��
2{՟�����0�a���aˁ*�3�I�3o�h7?�]��;���4恕�u���0Bk���w��:���r6�;�B�
D�i�C�؁ΐ5>OP�&Mk�M��#��X�7nsa~���Ӭp��xg�(�B�3�_��~x�ճ�o���x��S��V���TI�E���(;��=!��# �޼��ic�yc���-��V��3X9AC<�hC��CȦ~y�o'×���h2�0�!VX$)\�>t��i=�Loe�-��������2,AB�u�CEr6�)t� ��/*l7)!��;��u��'w�-���iهj�� �Ҵ�~X8.G-ԂJ��f�[ �|�C�vb��?gh��v��m#���~C�5#̇�l����Y���S�JRk)�%b_:�9��A�7�ݴ@03v�)(�b~n�t�g��a-.�%��N�kpi�|��/�m=���X��u֐F�'���LԻ��tPt�)|4J�i�Ye�#�����v$�;��1�F�3*�l@��#?$Q�7���>�Ƥ����ڒ�$6�3�}� �rʮD ��ȫ	����еp��_k@��i��pP�o��y)ke��Yj���z��1t��a�����
%�±�C����Li����VpQ��v@f�~���Ա�}�A1�"wA�m��(VS��Qs�t?R�-��:q�*^� ]��$AA�AG�H�҂|�'��@1�d�iP�z�'���$90���C�;#� �٩��'jJ�\�%\	k�R�����%�.:���C�&a� g�X�nC����Q��%>/g�My"ǫ{��-�n�{!p��3�6��-��z/�۱���1�N����/�3�^��d*^V���� Y���I:k6�T*y���c�\Ui�>�M�v_n�iMd�xL�o�
�h���T�@a��jxH�Dڙ�t1��O���'ۖ�U��6�n�����s���BB��ẻ���7ƃ) ��L�f�����E����A�))Wy�pK}L,��nK�H�r�_I
ъV�c�>���>�����T�ؘ��4���[�%��0�%M �oL�
���V��i�BS�� ��]!8+�9)꿼]�#U�����%7��~/ ��~L�+��C�4���߼����:��> ߍ����/ݔڲ�[&Q���>��|ǣ�p�A^Dw�֏��5�[��L,)܈��Ϛ�]�;��Nyo[~e����S�x0/wt̀}}!���-�����[�{����v�R�zu(�e����b,��Y�u'���/s4�%����<=����}�z����d���}�~S� #��q���.kaaZ��@�Ô�f��>i�6�קm���G9ЃJ��h�T����@��?�IN�
��j�w:kU��D��g)W�y����/JɘA_��m5 �[a��E���֋���1/6�ۦ���l|�����O�pd6	ۘ���gʲK�w��BM�a'Ö�@ց�vyn�*��Z/��g	ȼ��%�z �EF]��x5�����6\���UH/k{���b��Fl1,�뿴Ÿ��������K����0����L��� OY���V�8�&)��~_�Y��r6�ۅU٬�;G����Z��3�iIsM�])Ya����"DɃƮ�DB�#F�lu�������*8Ͷ�����
�zM|/v/g�@X��ŖR촁2�����}iV���a���P�wE�
����x��P�<�<nƂ��3l�NU�� ��u��\Q��~���d��B��{�%�Pd~�� ��ϭ$�fL�m�/��+C�fc��Na��E+�����9�	oG��3��>e~�23�/V-�72w�M�۟=���G\��;i��V��
�sX��d�o�,��?�۸�w���r�j��bϥ�M�?�8'�kԀ˕<j�>Z�+<�}J�R���u�u�`*�6�B3���&� #dk�5����6��Gc�W,�`#^(jx�cќe[l�&�v6�/�0X*>&����m��m�
�`!�%p�&PfT�Ɖ�(V �Fa��bc���@(�sv|�fK8�ܮ���l�
a?��:��	��]����~���B�)4�a��3�D�8��_*~B��K�K�B0c�G�N=58�����Q*	Z��34�\�\�k��c�H�s|���<-_��9u���8K���ި��Vl��L������ �B�G`�av�g�Bf' 0�n�����?!}���6��)9�v�J����+�ض��&�����B�3���I�F�"���>0�b�G )!�0��&�l{�vd���Pp�}����BI$4ݍ��}/���Xb��p-VN��u�p�P�pP�������7�T9Kr�j��<C^=e`'^v�m	 ����u�����3J ��!	�&�^wP�0A��P��8���O�tC�D6��G==�k������xAKUs�ٹ7��Y�T�іL�æP���@O�IȜ�ty��9��ߒ���t8z!��{�cI�x��R���"��(�FN�@\XX����5���q���}A��٣�H�f歟�����|A�*�v?Xyf�q���m���/����ɂr?�p���\UK�U�6�����\B�ap�g�jXϘa�!=jAލ�\�r&>���:�[{�ϟ�x�QP���0�o5\֭�!^!nw���OO�ai�>��i����0��sZ̊��׳fB��=G�wʊ}E!��넢ž`h�M��K���K��i�/2˴/&�]�u�)�������i���j9�80r��J�@���1l�!笠t�	i��x��l�L3���,ԁ�xUT.\pfr�r1��:�q�;�����ك{v[�� ��V��*X�Ga$rו)S���2਴�s� �e­��=�Xo��]��E0� �-�nm��D��%)��yݙb�|�]���z*4��S���7��9�H팚�7�o{Z�Wh=������':���D�n��:�eN�������@h�H>�%��; � Sl�0��%.|�A�J�����3"	�:�»��Sv4oʸD�)m'H�.�<F��orB5*9���>�t���Q>R)�BA>��%�?��o�e?�E��CC%<�B����gL�o�}���: �(����	���8����*B`շn~@�C�?�b�.����E���З$��60w!Ѹ����'�r�bjKiE���$���P���fPa��|G~g��E(lv�ܥ�#}�+>Zq�n�w3�c�1/͝�\;�C����JC	�|n�v�nW3���9If�zY��OY��;��
��y:��@)l�-�e��4�9�w���?V�+��)s������-�ұ�<\��WQo�{k��k	3YK�pU�� ��Jb�j\)v��|�����h�g�6��]?ݨЦ�wK�]���P�Z"���ufUF��Y�#v%��� ��_Xb�u�N����h���k�t��=뤑Iϖ0ք�D:I޽Mၢ�|Z�M}3�����9��D"�L��)!��Z����-�q�/�����ׄ�r�cx��Lq�$���b@I�~���֏z������&8)�P���m�o}���i<�y����������]���@�;��w�E�?:��=�6Z�Ju�3N�/(����.�E~<�`٬��c��3!�Jg�YL��z��@ѭsYVw���n���2�M�p,4O�ۣ�?�>�:�fą�ط���I�U�K������^�ǡP��$d+�x7��A@vR�?��~��n)5j#��2 >��K�j���]�+���kY�m8�_Dv��[q�Y�����@�>ٜ�t�1�Z=�d�˚�/	_��n��nM��4�Of�s4I|��{>� ��Q�⢚6֌9=���^O�v7_zj�΂��"X���t1���U����H�\E�^�?��k%P{)u�:<��d��T��N-����qC*<��1���'\��ыX8�CF��xk��M�)���P-ݘ�G���: '��rh>K�)߬�a��q�D/NE�
��ΰ��y��sW&�;G�����]v����\���/�輍�:&z홻4��%"#�[�o+��(e{�'4� �"���jw�%Q�1g2	"�e����A��v�ciF��v�߉�
����1�јQ�`b#��	}/�%��[M� �g��t#�d殡7��_Dڅ�F�H�y�3��!��� u���+�+�-u<�%�7�����l����q���w}b��4��]�T�"�}bSU�U"���D��t��p��F��J�Bd|g��k95�n�BY�ِWsk�����1�+`[UJg�[;�_�!k�\S��Qa( ��0�z>{ܟ�l�0X�V����0\X�u�(�1���?gsZ�b�0����4E���ɢO�:��-�ѩ$lei8�
�� �����#���L7�U:+E�h?�dx�N���y+���KB���W�z�A������XV/��/N���S��=LB�s�u_�C�b�?�����*�U'�ӱe�D�D�V����\�k#P:?S�F@�!�aID�Vn8�����$r{��R��0ĩK�K�x�gΓ��X�Q�
��e$����Wᬖ-B�}H�Nl��B�.,�A�6��[2����AϏo�Q�3��j!~�3]��[���m�w�R[�\�0��o���l�+e@ԕ. �c��x�$��̽�����[�Ky;<�q����8z�c�"8����BKHT�YA '�)ez� �b�J���{I���	%�QH?���ͮ��TBx����PDm<EH��Y���׍����2����f�#�,��A��3�z��Y���떱�9��j�e��D	ۈ:ƒ���0�Vy�$�D��Am.B��V��u�y,�3&Fm6���=��:�m�.��S��S�7Et>A8W1h���@m�ʽy���b�@H�L����?8|	&�!T^uz�@#���A��G]Bnl9tIhi��#X�j�vsH�V �"�a��CZ0v��+�<B�L��ĚT���J5��;N���3<�n���3� ��v�A��p�[3R�b%�ٺ퀔�F������W;�~��,j�>r����~+4'gױw�EO��*J=*�l/`�Nx�L�!-�5���С~(7��&�Py���~�]}��/�^1P�"���kn%����h�{��C,��R\�(��d�Oo�Kx�~T�F��v�t���
���P?#>|[�P�^�
��>p>m�mAg�2ev֯��>
S�����|LJl�a�Q2�+p����� �: ���٢�;��r����>�E�Yq|��-��Z�?J���uqj��,�Y
ӏ&%���;�X.E�#�$���j�ă�	��,��篳_�m��!nV컽=3lS�w2b�k'h���tۉ�W�dl���gx%4O����"ݠRk��T��h�n1�x`0�5���-�4�}/fd/�j�m&�?�?�Ƙ��*�H��n(�12���2��B+��N
J-fq�=]�I��M���߃dw�!x��B~s��&.b��Z�fƍ�����z���<�<J-��2�f��7)�a��$��e@-^�DkǎUʀr�zc�S1���r &�0���Ц+#�Mϩ�ښ��_	�+z������O���eCW�Ev;G�@a�G���e�If��x�Qv�;��QItxѭ�����1 �xI􈚍5��3m�DP�A`�8�O��xe��`.�X�V���l�)jC���@��)uu�����B� ֽ�,J�.��j��Ԍ4�S�I~	�E0�b��kWG��+�zo�����#:V*@���2��$�W=�e�vD�4��4'̚.m8�)�F��cłK�S�qb��b>E�!u*-'�$��;v) �9�v�`�r�#��=�]����i�{M:S�P���yQIO�a �|��	��vgVŨ$ o�k�LVUXq[�	�]�o��}+u|����yF�%_d�&�1�'�Mx���_Y�cn��z���W�S9yGU��Z~�����nq�S�ҥ��3"�&�&{���hu��c��b5̙ �^��yR7�|���]J{a�)ߔ���n�KuZ��
���&F�}�:k"gLZ����"���|�-�X���F�.w�,�p���0�c���g��N�,��dg"�V,�;H�B��!	NK��a�0��P݊��rf�u�V�Ţ:N! z��?�&�������k�չ�l�dlRp�V QÁ���iST^�a�%U�
;8"�LhS:+´̙d�7 �,����� H%�c��[�����Y'~K�T镽��3Ч��\��lڧ���׏�'Qo�[�X�#we�s[��_�K^��M��a����n��M�r9�-�P݌�Wf�C� �&�?��nJXJV�O���)�V/h��^h�W�x����K�A�
��L�y�b�������%�#Z��ۮU�Nz�����oo�6�:J�;J�!4z��`ۣ�$���`�$���]�tUf�/��a}h�^I	��h!4��O�=K�>P�[)1b:�[��IЂD��v�ٛ��eq�=
��9���5��f�<ֆ�(���?u� �im�\}~�Y{H��n[��θ�*Zm0:e<EA� �+��Q����)ޢSy�/.����b��h�&�QC���s���C�Bd�����yX�iV�/D0>V�T򑟏�6��ML�ԂN�R#�lg�0	�����B���	��'+Tu���sve �#��L@d"�^y�m͌p���������Gf�_��i�Xퟐ*'��d�%�B���x�@���'Brjd���`����M{�Q9���A���j:!f,�l�n��j�.ù�ܐD�G2�4�\�u�i�kP9��?�����Snyާ�����g��LJX�j��o�)<���K���K~F�'(_Q˜6d��}�&�O�`�AF�����m��2~�A���]4$��W2�C��"ji�k������e^a�L;���/4h(v�U ��[nڝ3JS˧�9�4�X�<;LjqG��2K+ɡ�@^��:�pV~ڑ裦!���������M1��g��~�a��#���q:��K��wB�VNMfH�,�_��W#�۫�S�Y)$���":�25��j�@c�,�[J�L����%� 9��yOӃ��7�H�JU�K�R F�_W#ǏU����Hyi�:�g~��+M)5UD���4��B*������h˓�2���7�(�k�/�7ñ�cwR�u��������7���RZ2�$��d7��mF����h+#b��N��2�ߐ�W��N�H&�no>�.�@�'�w� �&��_KX�iC�g�C
>D�^�p���Ec���ȣf���m?�bb�I_l 풱��8L=�z���d.w G�0�(k��Xނ0�I����g'��|�?�r���8�_�},c<s@��������ㅪb��UKu��H.b]Ibk԰W.��p�zP�2C;hS[8���?z����R��νk{!Z���2�+�5����i�5%�C��Eq,8x�����7'V�	�A��rd���!Z�k�_0G�P����$�eʻ.�N���k���My�8��)���d ���C[|7Aߧ��̜�I�z��
��?����I�]-���DM9+���/ܵ��1MNbjJ����i+B\E��M%Z�h�Ka��dU�O��2:{���M�&���������,+�	���<n��m��1�v`�Hw���g�_��I�'�-�^</��O[ǥL�����Q��F�^|M;��.A@��,���:�%N��/`�0?���J"-�v�FXpH8���:C��T���"���9�.��&�lb��	��7�C���D{�6Y&3�lЈ?�0���U���;T?j�r*_���=؇��@���L���m�Ka�?*��:w���g���#�2�Y����ꮩ_��7K�>FY<VsJ�V���?����RHW��>6D�X��~������AKa�~�,��k�RV��;�`�+KE	f�|8�r6pt��-V���.�n'�m�.9n��)7K����Ͷ��y<��Ʉ==M�����reN�;9��LP'}�E�:��jF�@M�hnV�<q��Ӥ��lZÄA~���<U�Ã�����&�:
E�K���3C~@m"��7q^�-���5Յ���c�6Aj]=K��Ю��[�{Ӛ���OT4uD��LF���o����\���|�!7�4|fB�w���y�$���v׸� �Oz>��������p���z�>�֮�y�2`�P,��ԡ襓��7�t�z����r0�֖�s���/�ܨ�v��_��K0*W�]�m�v{�<��!��3B&���U\e��a0t ��~�X�{�c_1���|�����M�NtI���`�fL��s�5O�'�S}�&���Z� ��1Z��ˡ|�|����G��g�O�yr��=�2v�z>�-5}f\V%��ե+n;��+�oE@'Y�����.O�: ���:�5 &6kxz���<w����y�G��r��9.�T�����g�
�ٺ9���r�t����T����"��c���w���'�L͇{Oywc�k;���H��w��͞H���" �r�83tY#�ȴ�`O�Ν�u&�:$����d���͒i�JՎ�y���B��\�TOLq +���j㛽/�'ЋM��d�˫�W`�BG�}�JUE������<��?��e6����r�A�S�t�U�Ri|N�%m���+�
ku �T��$X��6BM?�P��p�]s\���p�]�a
�Bh��P�n��J=4�]�/�� �%I�γ�>WdjU+Oc�骍��1R�V���.a�i���d��ҹ0�Fu&Pl_(<-����/������_����<�S85�I◌�;ԕ2�w�'[�7wv�'nO)-!+#��OĎp�����DóA�?�����n�4S���Y=�n��J�w�|��Z�����S�k�V�#��Yf�����)�f��YSDSk!Ԡ���h������v+X��o�'�.�_b2�At�</����t�m�L��m,��9���GS��&���/� !W:#tI��`nr�$�Y��f��p��)�dqݼ�@d%3�����o�N��A �L���Y��3�B��Cw��Յ7��>!v;�"�ݒ쒍X�k�
̻�s�!�x��H�B���^$T>�����ϑL�\kK�d�d��$S5�ޱs�3}���d�\	�hq$�:��R%�=oF�5H����w��B�e����9m�l�����T�$���%��N�;���fq9q)���{��u��
�F�o�V�^�q3�R���h�ƴ�_�M�lcI:I���s��HT�RJ�uL��Ŀ�0v[U.��&@ޭ��1�o��:�|���:�B��IO�3�n�tU1��D���������ɣ�b}x�q���"�>�>T��EπF���S�
=�$����8R���a�q*=Ot�&��<��r6���/���VAp뜡��.�:]�' �yb\�	{ ��fY̩U�gW%�e�"E������T��8�ğ�
�J�F�✕�[(�p�J�񟹩��$�XRwj���R*����e�%z��4���&�}�g3U8U��=JG����G���I�% ���KoO'��=r�!qpRm,T 6	���i}�?A����$��-���6��A����ġ%F���{ԑ�%ƚI�I�)';5N�@	�k�[�I�'�\:y��A��dm�T�ᨎӕ�����Fb�}
�2�]���(L��jT�-)���i�y����k�]����SP@�ߴDEq�-x�Ӭi��� R��M�����]��|al&�̧����d�,6q���'"�*u�2�$񩇉�r��V!mK��c�D��^ی�rт��&����}&�i�|�֩ҹ P��%{��Q$R�%�5�:��u��e��7L���&hP�{������ٔȖ/%)F�����(��_����x�!�CgbyM;(3��f�����\�&phw�Rᐭ"N�bR͇�����Cy��k�2�d�����!�`�V Mu�9�A��bh�d�+�$��gĢ\�@<+] �(t9���q��:&�G.��9X������r|�f�PV�u������<��U��s�E�߽9�;_�QT��Vj2_Х��c�������������E�"D�u��{;I�M$�>�� I�T�q�z'Q4F>M i �(�|F�Rd��^��#']��Uѣ:wڛh���#�'i�[�g��8X֜��A�w�i�����U��L<����{��Q�K!6z%��3��F#W?�q