��/  �X;4AP!���(��AаU=(f����Pk������Ѐ��Zϝ��NG�ɭ������-hZ׳;w�2��+s��8B𐓳Ӓ��$�c�} ��+��]E�%9Ɓ��P���0��9Ư>H�[�a�2�~��l�c2��E-�IQ�,�-i�K,:剛����K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!����ıL	���dG׉:�v�&7^ș��+�W1���_� ��Paj�u5�����Q��ߝN!(�F�C�R�������O$�����W9��	-�KT8q'�J��ل�)�\��Κ	U����VM��'(n=y
�ܡ�T�h�"@=֔�/q����=w�K5�@�ǻ�U�̅�/���1�I��P���D��!��]�1c��V�����4 Y��6�rrF�Ex���F�TT���&6l�'�c��~�ɞ�	��S��E���v��
s|gU�dG��7����d=y�]�D�h�/���a�2*���l��r$���9�vta��@3�!�Q��Nl����4J����{^"�{0IQb���̽���T�S̡c�r�5sޞ��x����B���d��S௒"�Ko͞����U������@�<|��a��
���PV�y��B
׸J0G� v��ʗ1�������H������'����<��)���H^��G�Nll�L����b�Β1�d*|��s��":'�I�R����?�M[��߮mě�Ƅ8=�H�>�r�.@=*�ɨd���)��5<̛�؆&��B¿$(�_.�����,z��}!����CU9�rL�A��N� ϝ��kt�9��, �	�9���%X�DK��Xt9ON�\�?��t��&�*e5R҅�����@�H�$��]Wg��w1���|� �ۓ%�#���PW:,��w��@9�,�ҷ������L�%i��Er�������4�ɶZ��,d�����hb�}� 1YY;���9xt�W}�걂��YYd��4����2�I!!s\���A����k	Q~ڴG)�L�M��bz�bǭ�����4;u �E�j��Np�r�[�ѧR�X%�A�R���0������>�|���v5��RE0` D�1��ay�ս�8����#ew �r�m��ܖ{���$]cb۱Ue�X�) ��qͥI�Q���6'�&��\^b�jqXחZ���N��!��H>�;��!�n���f��q>����ڤЌ`��Bt)p�"�:'Y�H�v��5�"��s93VϫY��GY��GA�c��S߿2dBVg�J��]�#�t9�ni�\�-k��	����HK�����-�'-�����t�k��8���\1���S�V&20ߙ ��E����B���r����,%�����ݮۦ��>T�j�P�R\�5p��IԌ'�R��7��W�����R>&��\� 1ߓ��Ned&��[a�#�j�����?������Yír�=�T+t>�CA�h�ן�[��b�g:ɴ��H�b�-����'�@Ϲ��G��rb6���K$Y^�. ����W�[JDmm�N8���Օ�����<uK�)6�IG�Xv�����[�~���GzY��b�j�v!/�������6�e��"!Xc�~�b��EcH��`�Ge�73ޯ8�G>���&��h:�<F�+�fc�(�����6���r��5?Q	����ӂ~>!Ͷ��� 9������tx�t�ޔ�4��Y��F����n� a������K���v�CW�=NH*�H{��W���:�qC"��zN%	_�K��y'�-;��|���&���ck�BX#ڔ8}J �^*�`O]�Yxf�s���\X���]�Х������գ����T+=�!M^}�89���{b�UVp:������ȣ�P��A����������