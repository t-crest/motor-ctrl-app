��/  h$�p�̦W���֫�hO�\S��F[P���!P�a}8�md:3��jc�M��F�������^t��3�%΁ �Mg��x�Q���w���|3��+Z��b���XP5��l�<љ�
azP&V{7ұ뛇A����R ~�wH̬�_<�8���~���š�K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<p�at*;%%���g�N�"���|�����Gw�+��݆(���7XmnA�=��o&#�]�z�5��;���oc�2�:�[�����;OP���yF<*��D��"��C�{�Ɠ@������o�Z;�j@�@ +�����`:�&s�G��}̷��Ǜjx*�&|rW��_t�*�-��⭣F@c�c�S���l�i���l���dC^h�w~��x	/����,Vo2U"q���Z5�U�ۂa]�Vܜ�t��dA�%�"q0,G|;�y�)tW!��qW�]�7����)��������L&��SE�V�-�&�zR���)A���-����˞Z��T����4��f�I8d�G�{`�N�-7�_��E�)�%���yZ#��c�������Tb@1
�V�T�Pt�ǈq�cP7|�&����<rU|��/�Sr^SRS��d�Z�jߪ)�3�.F	�0�[����#���q�D����幡�%�6�d��DV監4T�V �4}`�i���,�h��=�J=6G��ۂIRtWe3sO����X�;h����R�c����S�J�+lQ�K-(�ea�`@�����x��G�j�E�c���8�V�r�jDPҐ/�Ȋ�s���Fwo��%����״�������NH��*��ǎY�{᜵����م��L��jk޲?�y�'CǬ-M�T����vvZ�ۨH��h���澓��2����~�n<���3�0�����Ϣ,��|Lx��:���8^B�{b	�(����ս��Ь��*�a@�d��h�K���l�1i�������~��D!��.����w�������!3�qQ�*�0><r�C��k:��
.��Eot��T����b8��j�4��YP��b�ɚ6�<��%.v�ִ.4��X~�>ޝ��M��ΫF��l��X
G3���S`�jo�ȦKg�<�ʪ�R^u������:I�x�C�6��u�ڞ��}Ux%F�v���S�g����r��6�2n�i����3�fxP�T-����\�vr�Q�n����t?�r|Y�E�2��>���IQ��n�%�Ь[5�֚|#L�l��c�'�q8�d��Z]5�����M������S�����,���Yh��( �Y^���6��W[#D#��ONk��yRR�R��Ё�w��SN��P�.�)�ٛ�D��f�=Y�S�=�ò/���9<�=`� �zy�ϰ�R��\�ʻeVͻ�^���gB��.�] ���^��,��E��B���Z�"�Lg:/�er��YP��憬�.�rs�YQ�f�R���[����_���� N�ȯ�\�t�x�]�"Q
4�E�^;K�md�;U:�n0B��gK�{!_g,���[��(�tnVry;�'2ֵ�5�P����(�pe��Q̹TZ|]	>�U4�oҧ�f}ٓ7Z�᜶��	�®-2.���BR����K����r��V��-O�Ӓ6W*'x�A��{je�&����^p$��ؐO:ܫ�^m��9mH��%DH�ِ/b�������P��
�9���Y��@�PW:|��W��3;F-�(��K(�N�NbsO��5(�G��%ف+��n�)1�ڜ�m�8��/k��"CZ]!v�
y� ,%��P��h�Q|��S�w��4d$U����b�����j�v�Z��( �J�n���;�fjY$���sa�E���֡4��Xy� 2	�	"j{��ǟcN�e[�z����1�2�h����n�#��O�1~{�u���|g"��zi[߈_5yq� 
��fUrٔb/�C�j��^źOC����/ �D���5�)�L�T��B�p`�#�$s�b�jl�pP�[ˎ2,#1�|[y�ע��/�X&�
�#pg�x��I=��c2����5:�	��O�L{�X\b	���צ!q��k����(�~ށ
��PBy.Sg���8��UNM�(dK���࡭AC)9�<Ly����NZ�R�s�(�r+QC�Bm�t��~w�&��@@4wl�������.E��G��VWcW��~���h��d}yc�mA��l��T���St8��J�Ud�M�6�+�B!/Hb�����4��y8y%�H�n5q��2a:8w)�RE�+�Y�l��w���;����*~�3=��X9�زC&xV��[�x�Hn,�~�.�X��;�nrQ�Y��6}!��%��05'}�!�EqL��k.y
ؙ�@��1T�p�s� #A���eů����L<j�>XM�9y|[�ܹ��cV��7�Z�E��fۑx�ḱ�'���h�-��qMmf�?��1���U���Kl��F��D�}�JY��W����'�7�*������!�S���_C��n�_��M�VŶ��1Z�w��bP&i����@*0F������:�ugRZڨ��3ۏ,F���{G|�\F�+NC�H����HUh=`i��a1�9󆵺��7�"�wY?��n��aL20�R�����}�rsG�j'x�΢(�S�p��'v/l*��R�:AM���5�@Q~#g�}�����S(@�'�/h�nj�����݀���l���%�W�V{}����u�{��Z���8�Z�#��נQ��4o�/��
�������Qyqx(Mj�1#K�XJ1�۬���Ψ���.�����&I��Ss��Z���H���~��q��	�0k�����q�_�vE��v���c�C��ȓ�r���p����B�����[I�{Ϯ /��@V
c$c���i��$A�����/�))q`sJ� q�Ƥ��44c&����X,�P+��"&>0،��c�I�Af#jT���$RU�t4�QX�Ӵ��8�:��Au��sJ�Kh���S���Ռ+����V���t.ӟ��R��p�õb�|c��������Q)+fe���|`����xݠ�y�����8�}���*��N=��c-��ΉI�@,�>�K���m�;�����'��j��c ���IT��/i$��Ug�nE�s?��U��&�M��9�T�g�v�KO�����:˰_�<��V��Vx�B�����aIeX�W�|����Hj�I�<�a�.F�A�
�#�h��3����}�Z�o+����n�f"|�f>f�\M'��c2ִ@��~|��n�'W��{��faPGڇj�r����G�bs�;|!�-�jv�rE��P6Y�@d�m
�F�6��9��Dm���rZ�@���f�{T��%&�K�Υ��D��I=3n\��t��O�/��"�`�w�9
!l��T#��0�N�\eM�4��D��6��YW���ci���@R�}���
�~���n�6�tR������Nדnw�|L�|��P#�e���7�(�fO�U���Q�_O�dNS����IV9����};-�~S�v�>
��������I�1)��Na=�\��,�!%ʣB�1�9�G0C�n�������4
�K��֕�u�(�ᚯ���;���L3�(�/IO����(���0uÙ͂��F4,U"�3�dEN���b�z��
1c��Lgڳߊ���KuwiL������}_?���J�Y]�H���t2�>��K�
I=�QJ٩�;�1䇁�;���#���7b��T���I"�q�M�xY; �2������_nS���O��zy�(�,as+�v>�N6��E��*�^ʦ��PV�E�G��D���;~)�V8g�lk����V�����?y��xX��I��x��vr���Q�9(�FK?�j9��\]3׻vd�0��x�ǩCM�U�5�&sC�m�*�/ ��͖$9�ac?\(��$`�%y{Q�C��S���I���@�q�2���ul�E�?س��2�0�)&���;�V�`�!/�(;�
�N\���UO�d�;e��S�ALR�!"GƠܤǜ���]ޢ������mx���Z�\�u�P���E�Ty�����X��.h�j���Lb�p"CD�>���.�?o�������M�78���������
[�!�9u�]�wQ�'��A!]z����]R��3d<�G����h:��+5��>_�8*����;ί�����j�n 9?�L2�?|��::6�ch����FD1?�G���ʝ��ZkY/2Ӯ]V	C�B�- ��S�^��t�d�ނ�K����;6%�g�|�л2U�z�	��[�q��Q�U�?W�10�v���됞��(UH���G�1i�|��Q/�{��|]z�(}Pj4�7����%A�.�X�U1��/����,Y0�B�uL�al�EFKnHLi��������@9P|�o.�Y�&�6<-ќ=u�1��dWس�	����¹�B&��dTl�)���������~��aUS�Y�����#L>v�C�i�|����^.��c�z$YC���폿�H�����|_zG���D%���L�bi��6<&%��@�:�ӧ��$a��S�­��QO�a���7���������)����a��e�ne���WRN�D�WT2���i4L����۲�êjC9������O��9�yI�Dʯ�;�'?�$�l'��2r+�#q��_P,��B�[���=Ñ������o4�v>ZB'���� �;o��M4ᚠ�GN��84T6��g��1��;��}UF=��&qFL:���}l����vjРj�2		�0���WBPƕT��-S�F��X#b�����|����rx�\�{P�\�8`���^�D�S�d/�����1ͧ�n��E�x�&�1��G�=��ˣ���|x�Nmw��-�;��X������)忣t�M�#��V��u��w�C�Π$-��v��v@��:h!�W[f�-��z`���\�\����v�8a��,��n=~Wn�]��y��R�viȖ0#��L���<�b��=�;H)_�p��Yw m��鱕���(t�0"�J�i*p�N�G���H9���^��R���T9�p���;���A�pk���X�H�3
��I�1>jQ0`jq�i�$u�b����+)�nm������TJ�O�s��,O�J���I��+`���"������C@!
��B_�Q��
(��i�/9^��]b�Z�X���cH��9��Zv�9����>���"��M�p�mI��i�Y1��upFp89������N6+w�e��D�c2�}�"��W ����5f_���jk��3���a�x��T)^xK��Q��L#~�ׂ:T�y]�`���μ��ČO�%˃hfD��L��0�bڑ|����� �T9FO�^�j�U^��܂~��1~l3�Q�7W�U�qU�[��:�?��jP��ȭ��z���t����_y:�Un�i<Bq�<�v�<�3~Ӑ������<l���x�/*�	��23[3 �=���2�B���W�˼|��h� �1��ƫ���#�^�6U�gIS3���2��]��N��4�w�	����"p�ʎ˺�c�(�,"G���㘁)ڼ�c�qNi>�3O�"����ez�$�P��c2E���G���U�	l�T��qd�c�n3B��UŁ3��U`E��VIa���:@2�%g�`��2�+7)��Z��4��IȜ�Pt��-��i�ι��CL�dAdXaUޏؓ�-^
�k�W���&���\H�/�.u���5��@�H���4Vw��L|��TH�?$i�u�0.�$�fR*�ҵ���+e-YX�M����}0i9 �V��������_�N��PV���훡� ����?�pd[�cK ԏ��j\FE#��a��ą}i_�HM%Mr#c�������ƦA���`-���i��lyp&����6BPv�-_p�H��9��A�%<�O]]�"�Ҹ��õ>T���>�=���Be�F�do��� ������%�[bۜ[��w��0qbi4WU hBH����=�(���cH��$ъN?m��4O��%A�(�Se�uͪs�^�b��^���֮��`b��-@*V��-lVDxu N�����U��V�M�Γe��~�������f�j��٘hL�/^��4��~�6Z�������TW���?fRkE���ak}*�S:���/�����9��Q�-��<<Y<�e7�@ε!>�s�ǩ{'�F/�l��@si��3/�#2"��n;�:!g�*ի�<'g��=��	�C��6s�rR@�N��>q~�>ݣך�1E%C$�ܴ�SB��/$�f$V�f�a��R��,Z�M�&�H lg.?n�(����-]2�5ga���<Ay�>[��A;��p����&U�q^,)��FD�c��eEjBiu	ʄ��'�O9Z}OH�
�����%�>$S���Y-�}��USWog�²e��zD�_Q%}�]@���eD�-�Z����w` ��[��Ԇc ��j�Fg[��+x��p�D1��|��a7R��gG�4S�ˉ~&��ڟ�����'`+�T�4���ݞ���"2���J�f	AoE�=�A�#c�z.n�1��eP}Ha�x�Jݟ�⼁cֱ�`��Ke�L����̄Q2R1�(�*�=(��X,ƌӵ�"�VZ�ki��� �ؗA@�v�,����Q�b��Q���^��R�b<������|2x��5l��%� ;ބ��3N	�|�mq�ۜ �x�Z�H�c��
��X??=ӡ=�h`�FPj�����C��1�o�a��i�C�$�w�N�hW�?�Z�~aJ=��Ql��8��.�n�J�����L���B�iq�J0��k�30�ڛa
������M�Md�C�/E{���-�:D�B:Đ�H  ����@$�s�b�S9����1}�:�������S%�0�ݬƐZo����,�S�ܿ$ay�r\�Y��1X>g�Xy���|ps6$(�1w ��x���5!gx_§�aZ�)�P�����io�����R7Sl�O��b������L�~�I\�Sğ�Q�/{P�/1��3�
<�����*Pl�'�Pe�C���F<����nc�@�0�X����������������T��0ة�J`@/��&?�0(>G��k.��!��A{��I�Imr��M����X�Ӻ�eUGkq1P��G����4 8��	
N�
j��mnr�P���1�5�o�s��E�f~ƬSbB�@?�D�G�F�Z���y�Z4ۏ��lט\��U63�ĮN�����$�� ��H�Jd8��p�oc�~�T����1����'�k��_)����R���кbv����!!��r�#�넜o٦
S?P*��9��擣��� _}���{Cs��r\��J8�<S�5
���˞��O����"��fߔtO˂p�.�TW�@�����up�؞��̉uR�{�,
�J�8FǷ�_��|���u;��� ˗~6�5�� �����6�[cx<�cw�#W:L0W3\)��O�j�h��� �/V���J��F��7��ر�����an
H9�h���Bl��Д�3@�� �S��&F���9K�Q�֮�D��_&3�#�h���nÒ��_6�����_Ѷ���aM������D5J�v�{q6E�7��g}ߤ�n�4f���
Q��j}C'%.t�uS}�<�(]��|A�����!�W�h�z�W�,;��ຬ��.��=̍d��V?�3\mpb~�#�(�y/$���ʽ\ 0i��<�0#�����!���Uʀ/ bU� 1�G�%�E�lTS��Ⓕ�)��	�>�t��!�4Zc
�Td���4��8b�4�f$�
�'7������P�J��ů�X��'!��k�y���9Nt��%C}�!8,��Nv��Z���ֲH���@�u//QF �	�7�~�D4��e_¦2�ol���D�.�89ȏ��@��FJ��"��VT\���oq@���M���֑D"Wx:b�S#k��W����J���b��
�\	{"�%A�@�-��Ԧ�>�{�{�5@)�B��7���_��9 �A�8�}�tv)[��p�ױ�l�\�!�5��!����{X�\�4�����%/y�2��u��������u���$,f�zl��'�e�71�ގ?#.���v�(��5A�Un�ɼ;H�7&���{�4m�G���߈ �(�m,���	p�%,|�e��K�/h�^$��ĥ����泹9pe"z8�o����y�B�Ŀ�_���sò�|�|�G�&�j%��a�&������Y���'P"��!]�G���W�P8Bm��dytE������jU�����#�^rNU�Y[Y�&=�O�W�Q)�b��o}�MuT��Q�
��Nc�T���C%{r�/y��N�������Qj��N d������8�6������!�n�ièN�[K���)��x����%��L���^��_KQS�ŕ7.D���4Q���4j�3[\���U]E��1Mн񪬎��Ȳ}��5�~e��?O0���b|� ����<?a���#�Ѱ�R�/�c�_��O�N��h0�xg��x4{�5y����gUdG��'�R	u��?�FStj4�r-
G]덴b����+U}r�:�Y	��z���"�Ǟ�̭[�j��8]��I�Rj�/�`�f�����S�!@(V�����кz�f,��6�����@�(�t�U��Ȍ8 S_�u���y�w���0D��j�j��.�����Y# @�Ǎ�5L�pi�F���N���C�}���Y���@%]�	y/X&�~�ț�3��Ğ�aF�)Cmp�۰��5"?�Q�ݡ��?fӥ
�3�.�/�مd|�0�,����`	�`��/�el����+[�
�qܙ?0�q^l��M��@k�}@M��j_�0�kg��9ص��8a���]�<�fC��Y.zV����Y�?����`2�����-��P���27� ��St���i����!?��!z�N�2�z�,�$�&d[7�� n�r���S-n$��͂]�-��RN3�e���`��B�Z{^���/n�WT�#{��"&�r�7��d(�EI笔!�oM��xzG�����d�M3��)0��;��DG�u|hXqe���*;�;b�[�xe���0��il݉N4�f�]i5�e4F��Cؓz�E�������J�Y�����zXM��`ݞ<����/,�IWAs�3rG��~d�����OE��AH��/��Z�۴��a*��!p�z�_��L�y�6�SQ���o�Y`��L	-���n�(�F��=��u5���(LOIML[09#����3�!g�c���r�*�=dq�(^N"$
l6}@[[��U����X��vE��m�x'�U��Y�$�2�qɪ��(n�U9���е�.s��&ifĤz�Eq�f'�V�z�.s�8��E��=�jC��}X���Y��^�C���;�R?h9���H\1��rKE�S�N��z�j`�/paMg���u:9��r��n��I7HI���(\V����j�ݟL���4N��;%��WR��X� (2j@� �N&��=�s�7��ܪ��7�v?Ȩ�e�TK@h���&���xu(��P$c`���Tci����dy���ن�yR췥un���ҶӨ��1k�Ez�`h�iK�M�������5����ڦT/{ka��u���#+J�l�k�JƤ.�,��S�{S����p����l��>�郊�I&���{	�W�&�$݅�n�%%��+���/WʐoR�Y��ݓ4����r5�P~LA��%�j�|��ݦu~��F7�μ���BZP=#n忞�Y&rQ]m�-`~5&�)�	ͷ&�`9��jS?|A�0�z�>�,���e�a �&�h�Y@u
O�wo.�6�`d��V��cƥ\�Hh�z~ђo
iCP�D�P�9�e�vZV�,�"���o�t#w��U�m��$�f�R7��)X#��1�$�A��}�^l�s�p3� n�x|�����tr_������`|�Ĉ�NG,Q���ӄe���[O��W��<�T�W���ǔUty����^�&�o׀��+1���0�����'ܷ��4Y������;���T�Юk��}�*�4Ђ鿒�<0x�2N�_I�C�l��ݶ,T�T`o�Z�pi��xR,�
X^	�g=�S�u�#�+�)��6T��闯���w� ���fE�����2F�٬�TF��")�yּw��;�i�w��X:	���;���_��A6b��=�q�t���Ch������TD�&�b1 ������5���v����]؉���U��s�Ҏ�CU;q\-xq�}�ɖK�ӏpS�� o�����?6mj(��F!�:��hs�;��P���H2S�`H��9��|�<�#W�mr�n�^�x�wD,;QK��O>�Sv?�M>�x���ӂ��P�l��qMR��a��E�ܒAq�N��g��צ46(�8�4{b�M�ҟ�橗L���]ܐ!8��8�8���=�_���`m8���ʁ���~pZxk�>�oV����E"��o���%�(��T�h&�����o� 氺��e���R��4b�ה32M�h>Y�ƌ���!�����@e��M�����Y��;��h�^>,��L;٤.��nbuo�Ң�x��3�0ZZ�1�tM��/�-�]�c���]�rX����E�\,�怛pM�5�r�.K7����/X2��v��'�)�d��'����dIw:�4R��?B=�2����5V�;���g�X�m�ƾ�;:Tp��O5t18賞MT�(OPalc~�?\�+��p-�%�[�:�Ě��s㺟�^�=ֱ���U5j�3?���_
q�0�=�m^B.�\\�ly^%����n{�����:@(�3q�Ƌ^쁒~��:���%���K%�h�"���5F�ҩ�K������3XIB��+ڱ|�$6�Ņ�cY 'O� &�-mw�So�l<�{�����Ճ�h��I����>.\[	|uqL��#X�r��uII;��Q�y@~�#�>��8z�K��^��4�����=�o�2�[�����$U-��krMx���i��:�"m7�>�!�&��h�������Hi�X���[���R̢�K�<�G"��w���9�䄠�_u8+
~�ޙ��p�z�a��O�|�eW��թ�a6�j��iւ����3��-tl\\�}���������E�wϧl��G� �U�! ��sliedjR��N%5�OT�n���n��k^��J�d(���;��j��y���:Uz/Ǖ����(��� �$��{Z��`��Z��n�G�?�E�pBi�A����!H����̀�/=`�b	a'j#�n5�oTп��fb�1n�b���
Cpm�LL�kp�wFH��7�{�4�҇�d��atp��r��+ʜ�����D%��!�u&7f'V������(~��5o$%���\�#�Ì�_���*���!�g����mܯEq1�*��7�B�����3TJGC���ǸI�N�L���4�� i#H����W��D7X�!6����Y���瑀u{-�n�*��S�$?��R�i<tT��U�3׎姢�}+��G�o��(7
�q�T����Hܴ&Z�?�h�����1=����x��)}TI�F�]��+���}+vVg>�;�o�og�j~W%���Ya�|��㟿��c(����A�*��~�QCJ������!�Y'�6@l�!,@�{�ӊ��@�.���TV{��Uָ�7ľ.�`��%q�t����K��Ikԣ����Y2Z��Д�K��qж�Vה �Q�ƽ�{�8ΰ�g��z��9��%ďvI��?�T5�� �?{LR�m�q�v"|�*'^cD�UJTa�ח�ʴl��VA
��^�����lC�k����g�n���S� �Č_q~(�`�j��#��{ g�� ���y�!��_q�n�I���aI "Y0rj���>����DWq�q�hJ���N�j!`ڴ�|��3��|�[�X� ;p���Ʉ��g�X6o��%��Ů��]OB0���m�2d�q�4G�y�d��Q�������m��|�x�X��]�t�.Uh�̽��ܕ�D��a�\
���H!����2�$M������	4�6� ݍCߏ�hM�����%��"
���[����&�n����֦��8㒟�,}9��R��(B�o&�.���~�*�5�G����eCg=8�k�y�քLh����X5?�!�A����d�jƗ��?l�jl���K��@�3i�G�Z��40� �k$Xp`\�O(q	�ł����[��81��2�����&m���؁�"M���
к�����p�/5j ߺP�t��0	l�:%�l�w�Q�t*�B�]b˼7��T�r���`�;�E5�f�M|	�+�ޑ�ƨʼӠ��]�t�cK�_��Ǣذ� �^����i,69�����>�p���\�~+3��8?���<�sܛW�=sj=#�К^_������A�%����l9���9�h8'5��͙�m�(M��S�Xe,(�e� 1�![��ph�3�&@x�s7��`�	�������7Q~и��8�ӗ�V�Rx�(Y<|p�w�O;8��1�s��d�G�y��I��w'���2�E,"̱/��f�S����Y���j���؈PCٔ��3��Z��G t�x?1W�9�H�#6��t��3��/x+�2�%L^��	�C�q<$�K���9�Q�'�k���	5V�4���)JAy\�G$X; ���q��oϛ� ��=��0�������ZC�aʕެ�*rb ����o�ǈC	�9sۊ\B���耈�N����<O��>~�3HC�K���M�Ρ��FQ��2�kۜ�&�ܗ�d	Ï:�0q�dɈVF3���f헸�/{z��Y�E���!�Fd��0��\�Λ����*��A��A����K��V�i��<�)@1�D����/×��e��� �>G��9Q��AN�H�#��u/m���H?Z ������r������D�~�w��cʻ�ث�v?
ꯛ��n9x�lv$�#k��kL(��.����4��K!y�w'��d�u&�F����0�;����ad�,7-s'�
ťyب��
å?Ȍ�3��q�n<��-�Ag�(ח |��j�٥�����'��W9� $˶V��t�g�����	9��{�e�҄�D;e��M^�9�(Dx*���R��� �ES9���j�4G�.�ysf�/\� sq*���i��bͰ�6�+ʏ�����)e7`gbNa^��a��o�M���xɁe�����y;Y���Ap_�v
�[���/��,���r���$�S�!��:�/����ec�(݀�"*�4��ߣ�K.#l�/Ղ|p�i�w��OO�*U�u:ٮ�=8(�q���߽9��]����l��N�\��������Q.E�S�C������$/+g���f��'P�*|bӥ9L�iC��%���ﰺ���3�;`?5��
�Uh���q�`��Ȝ��y����BpT� ����Χ�W<����NHVY�|�|����ЧG�\��<�G1�� ����u��g�����O��{$�neC�Xe[�Һb葊T�e�Phc��L�r�m���e�V\����:L��VwP���+N�ʁΫ\�+���TXW�#���m�KH椢�+��u9�PM�6�/�=�������4�p٫��6�VO�XyAci�p����@�2U�ݽ}���rQ%4Bٮ�#I�Go@��Ϥ�-=uFצ�;���
�fN��{|��=t�>[:1��wԳ�zƵ%�St�S�������C��C�(�r�H+�/���s%ۿ�g�O��o]��h���Y�!s�E~��-������=�-JD��b�b���w<4 ���l��Ĝ
��2�� �8v�ׯ���q�i:�+��\��x��
-)�j�� @�"Y���qz]\���f<�"��ct�2���-���Rj����tI�����<g!5ph�}�����U����V��栾�v)�^#���E)@��H[}��o��0�#�yDE�oo��x�"M�2l[~�I'i��DK���L�1&���-(RJ��
]D�� Y��ɑ>�0�A����>Szs�\�ѭ�:H�����٣�-7v�7��!�
>����юl�ӃW���Xq� �&�=pG������71�4Ė�X��+�@DT~甾3"E�n;y����H�=�=���%�	���A���̆���ɵ����n��6H��߀ �[pe�}E�փ~$���\k��F�������*X�#�X�+�J���!�H���jF��Q�R8<���$%��<o	�`al��l�s��=��V�gc�:�-��oe�9��ؓ:�$F%�N��vh8-<�6�l]]����|
J��|fw7ú���"�-K�/GB"�d:���cZ	��=�*1���b,L}�X��7�\����~����9������V�1C̨{&��ȱ�zʽ9���3��@�4Vl<v�5�M�Be�:�z(�k���r��څ��5ރ���s��[E&g��c��yZ_7�8�m�h��1��ǥg�L#X_籧^��|'y�A�.`U���ZG�$@/A�Tܽ3���7�E$���/o��聁��V�����gd�ƠoMF_���� �Wn���߄�Y���\�=��mQb�T!ٚ!���e诘V�]1i��+5U��d8v�kT�}lm V�x�Xٜa]����j�~[A�U3ͧm�A�nk�f���&�˥���E�Q]=٢�f.�ۋ��	�̯��[�F��r�v���j�a8�_�lV�[���{����»���y�	�k���tlф����A��^�"s��C�p0$۰��ϰ5@cu[�nB	�S�ϊmQ_<�}�F�?�$!�P�����*DX ��	}�����u[Z7}~C� x@'���ee /#���;�
Y8��}"����bϊnT@k�J��v6�)�!Rk�(��K���X�hnq����?�TM!�%6*����I��\�)|�#�X�14ᦹP�|�nwN}��+�z��)t�@�v����à3�V0l����#}�7')qA�>I!���S�z��H�����H�s�##�Ј�N-���~'N��޺��17~	������ 6�8W*4Ju�'k�8zW�\�D�b��Pͫl�گ����G��́�Dƃ����!v�+a�n��x@�<�fZ!�@����q�~�(s'���,���oF	?{%�01KME uZ�[k[��u������e� 6U���E6b(� ���KݑG��V�KP�B���/ѭ�oc"�����SI�}�(�Rn��q�#R <qCS�I͒�?XX�e����4�	*!JM��!��(�/����8'!���֛�M�ΠZ�$@.���1�8�O|���"�������e%���.ޅ}���h&����@P'��L�E����7�������_���,��$	d��W�Fu�`n������c��bh��i^2`����bj#*�&a�û�F�_��Ӏ����@*aX}�#��B ��Q�����P���ҳݘJmZ����Ť����O������9���t�ri�p�3#�ni%��=�uw�h��R��,m8�I��|�^(0��R��8��w����2m굿�4-��r!���-�u^���*�ۇLe��S!}�������]_H�5��h��W!x&&�I�_ad��u�g(�u	��5�.�ӴH�|��S�*LCg�g��v3X�j��TY�n��=���^�� �)���S��c��Y��d�H��	v�u��)�m�zE׬����m3�	�P:�|� v퇊P|�h�nzx%0{�E����5�xY�ӛ;���P8����w�WE����7��7b,�o�&�9'=R����s���k�$��-�/�򖚊9�r����GjMο�?���߬������>k༻�́���[$�|�w���#Л,��k)���sv�o<�9𬏪�RA�/?��&4����؈Q�Ȁ�a�3�+i�?kg�T?!�	M�&X�I6M5���ߖ>���r�����q>�����'�|�_�\8���� ���]���0�5,����[��o���T�5MZ� �}Qt��
�i=�A��,�Sip>��C��dW�p�G(;��^�|��p���F���J�36��׀�u��$ؐ�D�ap���F������ɤi��'��3����<�Sv_��^���Ġ���H�R"_/Jȋ�I��K5z�6��A9�fhd�a���l��k[@����ǧVy����u���R���Ly��ɋf��>��3�4�A̰���W�Ê�"��@��!S&�����p4?Ǿ���#:"���un/i���X\�L�=m��д5�op{{��V�۔��ֲ��D��뢡c@"Z�r �'��5��"NHSDȡO�VIQ"�I��|����d�W0<	OQi���U���"!��GYL�u�� P_�g��:C�R�RVW4xn8��J	�3�5[��k%_���l��q�.�,
�q�(j4ƽ�}������E���~b�х���#	؁��{���o`���fD���ϫ�}�C4�V�"����WI��/��aY2���pb�s4˄O=��)'(�s�D�s͵#bf袴�3�� �6�龍����R�+D�h�S�ۢF,����$^�R�X��)8m󺞽*8=��� �D(#gVJ���MvǪR6�S���8�
�����h
K�W�D&���\����y�P���kS6�hA
w��Z�DrJ,V��ߤ1S@�Rr$�ޑ&'�r��c����X�UYD'쟫����7��RȌC���$��Wn���Q��*ҕ�R�'��ӝ���IO�C��G�}�yQƭ%�l0	¿��㧖 r�K"S��<@��xG釬T������f��S�5[��� �ϣ�M-�w^���f�V����C	n{+���=\+����8`@L[�0v,lzq��� �3@�68��$��k#m,&���uh�xW�j }��QK�N1s<��ê�R�c֪2�����l��<3\���Fϫ��,8�%W(<ʆ�ћKޕV�.b. �!g��i�~�,Ev�a)�=n��S���{���>A��Ē��J���YiuJRע��/ڎ�7�.�$Q��L��"���55���_�p��G9��8?-s�{��'�A�f���YK u�����\G������I0TRO���.5Uie[��v��&�pQ�i���]*�;�eu:
M@T�ކ��|~��-��I(\i#�&3���$��/;������\��::����/rm�oK`t�oJ��1袰��3������9�Ǡ�;}��!� ���"����r�������+��V��DW�J�;�p��4�ÌL,��dX���ᭇ����fD|�s��5	<���AS(���~\ ��?����fus�~����/�©���Ybĉ+d0cS����L1;Zwx��E<F]�~����o���*�.���18˿j�E��Rju|�E�w�ߟ����]\� ��X�/�J���v��Eżr�2D�5���p{Y�9�4�uC7폭���p���*�ѾVsgT�9 ͋�������!���7��'�M��l^y�Y���{�p�1Jpo��ooAM�^h�/4���ą��}�c}��8
�1����ƙ|���ah��#�b����Tcxs-M���,�"|
��Rj�cy�mY��;����MJf�E�snف�J�]$��{O���}�k�2!\~g�9�mOK�D||�I�|Z
t�zSd\7����)���]c̕�)y:����׫�4=�O���?{n��4O�̟�>;�lm�� ]�D�ټ؋��� ������͇������%"lehd���0���2�}�b5^j��Y����{��|�!87w_�G�N������-O_h��6|�:m����>x�P=��
_6�{�Rn������smR�W��|���֋�i��x����u�	m>�4.�'~,����-i�oI�<�ь��\����)�>M�W6�w��w�/��g2��hYp��8�	�  B�tnˍ��
c�;�[��.�|�yp�s{#�b254	�����yVw��hV+�;2����s�/�nH�D��)1z��Cx�g��|��4��nP���KE33n[3�|6b�v5�_�2�a�����%E+��};	�mߜ�j�N��mb��7x������r�9�ek�2��^$�k��9�`��uK��"�����.�vZ��}��^�ʍ���H��6�q���k��s������O.˗��&7��.�o���DIWY t{�-��[M�� I[6&t}&��	�°$��S��"���CV�����7�K����<c|�B!gTFƻ�������R�Qԛq����ܱ�S©Nb�M]�uI���<(Bԓ��{HT~��B$�R�?gڧ�p�:v��	JJaϸ��I��Nx�	y�;�:Z�޳���JP]��
M�1�O�e�H���
C�ڳn�u\�&����P_�#�v ,�R1�x+��n�߶���i�4�F���|�e�Z�q�w��эE�E�����U����E�={��Kq?J��2�g\�=��(�v5�����-W{JOXS�	�GRD'�A�E��Z3��ԯf���		��-։�5*���R"�zH8"©��څc0����'"�pE#<���џy�~�dټ�bTwð-l�ipo-Y��O}�.,0��H�� �_��W�q�IV�].i;�М�'ݼz}��yw/�U�؈�&o�q'���J� RCb��UK���0�{�V��>$G5��QK�|���Md[�
��Q"����6���ɬS�� �&*w"��\�=8���6�@�S�z�y>�|}����=�����5���Ob�	����(�O��I�����d������a�ޑj��}NRp�)mD�a���١��6�����Q��cm��	�9"���� <��G!g����tAY��guF�ff��O�Q
PX��������p^s)���{յ/Yu8P�J-����ع�{i]��� �n��{�j���m�EsbOӆ *�dT��9z&[b��w�-�|x*�)%bm���Tڟ��H�G\&g��&mDLk=k:uΎ�#l9X�9��hKU����������&00c �"�� �GN��c@�֜Ѩ`Tkm�J��o@z�O�D(�/��jޖF�w��ο�il�iқ�<�R��g�� ��%�j���tj�f{�K�h���x�����_��4@�L����0]��Hz~Y�@q�֑2�'�U�7혡Ԑ*uq[_)\��fKk��P��\\o�Y���Db�4��'.�#���������u{��>��]
�NX?��z=*�D��I�bk�$�[����v]Rw	�D2Ձf�B0i�����S�H����r�U?'�\(L��!�y��.�Q5�VJY �t�4�ކ��^:���A�Np��~��(!�Et�K� ��/���g՟�Ҟx}.�{�V�O�3�'g��ᔆ���Q�/�~hY�����9 ;�
�:��~.���"�J2k�GW_�W�$8�QӍt�ʶߣ���z�&E�*���F�=^؎ש���Z._��3'� ՛�`�NW��{xg[�6��a	&��]@�r$f(������Y,���?�������?5D>�	�I-��J��l$�vEc�s9��g�c�#`�������U]�
%?\�xJ �B�6ɿ�%lY�i���#[�й�:��m`�r;m�#����w;�m�g�����!�y�����(0n��c��jSN��"��m}�iF�0�N����/V}p�q4�ޫd���?�)�����bl-"e�o��&g�G�':U��o~�2�4~4mӽ�T6�BfMe\����G~uS�f��� �ϵ�<�A5=2����J�����2p:w��d�S�EӘ�LDQb�VM^%X�#�b(J�I5�)uv���(^��r�S�?e����/nR	-7�IG��~�3�j2�"_�Ф��WÇ?=
���4����J#���M�M�-�D�	3�2�ߖ�w�v�*�a��؟�=����O���n�`�{��/��Z�]b��n@�C��"���[+{���˘"��+HT��`�1���]���/�g3o~z�0#�it�4]{�^�-�N����F�o�{8X�P?&��C))ET�H��ω��M���o�!#61�oSz
�ai'Q+��b�>{�Gن�cvv6'�6]�a,�wqʤW���V}3��hE���D��6\��n�'����'���V���Vdw�i����`<h[Tiȭ������f�I̺�fq_8s��e<Y�y.b@�T���<Д�΁�49:��)�Ft�꧛

��	�d�)V�'�x>*���h��٘���M��5���ˇ��$.ʫ_n���a�:"n�)��S�J��l��9�4l�@n~� ��ۿ-� La��@E����ZЈ�:+���x5L��|�Wt�����Ң�K�+���_���/�UppK�pV�}.Ƕ�o����_H���pX�F�-a�U�*H�p�T�B�_s����逸�L�7�O�3p�Ξ>H�!88yh*E�62H��pul��sq/���L�Qr&��&n(��.vp'��R?�#����ΊB���1K@����;K#iY-��K�rz�ݾ�� ���j��������c�ā�π�35�T���9�Ҕh�8�w���
�U#R;����wˑ��^jA� ��d$�6S�����VJC�$��a?�Qr	T�?��\����$Р�o��aP�SiJ��]�p0���M��;�7��L�<h�8�]k_H���"	��߲	?2
g�A#�qD�L���˻^%�nŢ�������yO�1��z�8�O���"�˹f��ȓ�q
3�fa���r��+� � ����c�Og�M?�id>��3ΔJ��}_��]��/6d�j��;������>Y�#[������~Й�y��|��*_�~ ������Ȣ�':{/�$ޱ�{�,��������vz|[t�q����D龩�!�q�;�a�̜��;��S4m8x�����RqU�mM����w�h�������;Kj�7N6Q���n�o^�>uV؜aLΉ!/�������!�ϖ �300�\�WY��"�3����/�U�j"��w`�"����� �P4 $%B��v�a��Mq�Z�R�y��}��O9���Lcu��N�� l�k@�R�A瓤S��ܜ�ez��,��W��k���w�����O����a����[D�JQ����gq��6�i��-Ac�����r�!�k��g3d�L������5���T� +���	%r��fS��~?���� >Iv�w{�X\���8�?�����S��Ӡ꜆�ث	M�=	�/��.���4q8���.���|c�P�"�r;���B�Z~�OR��)�L�D�?T�V$Jm�c]��n?"_b�)�j�����#���G���ʶK���������M����Ƙ߫�tx��s]6�@,i����9��P�N����W���3I?��ۺjȌH~&E1���m�l�����S�6�M�� }�"��_�(4��N�O��МO���|a�8�c���WVCa�F�o\�%tJ��&M	��;QW��J	㕪(1#��S0��x�
bU��p�W�ԟ|�w�ۜ��漵�&�#pI�13�B~4��]���.]~xk��M_�c��jBpm��@YJrO��NZ�y���!�������1��9j뚒��2�A�D}LJf�O�E�<3J���L�j�(��o�>��U2#�WK= kd��;�	�wJR�<���. ����Y��9S��(�}]�B�N�/�|��=�ZQO��:o��h�Ţel+��:�iѿ��������*��/�L�����,y���~�}K}�2��E��5�
�>˻�\�����~*�g4�� ��-�`�����܋����2��M��>=�� z�k,�����ۛO����>S_�ה���A��h�^ �0Y��5\G(g/>[��E�\��=����8����J�ay��h��~�M��p$�M��6������u��f�Z$��WHxo���ּ������Z]~����(Հ���E����l�ǽ��6��i@Wb�|j��v\9�k�&R��
�̜*IC
M�Z�49d���}�,��	\�s]M+A�+ Q���|G�UF+_ۊG#��%���Q�\�0�9��MmFM� �AT�+�U��Fk�+�j�` '��1��&��/숉�R�	�]����S
��5����נ����(D'�i,?�3���1s{1*X]�:
`��CeԖ��br���F��C�'o�T�#dN�r`@���dǥe�*�:�)�C*�bK��{�x|����`��y���ˑ��3� уҭU.��H�'ԹXW��t,r��1����Ci��B�6�
�	P�)%�b��@_zB��ǝ3� �i�����u�����2�hW�;G1�(�KAH�>kǰw��"�Uz{	�r�C���s�7���U��n[�}��^�N�0��	`�U݇���zǬR*���fZAa�f�NO|n9�.��J�����P�9"�.�E�z�=�f��JK�$1[��2�˽'$���9��D�`[�3Róͺ��������L���>A�@`�u�t8W+��5ݣ�.���V����X�VJJ�3}�O@ߩ���c��9���ΰ�@�K^�?�]A����Mt#)Y$����3NM n>Z���if��E(_ۢ���< p��%�j9(j*;�i����)a7�ѩ��hJ�zNm<���V�8�CF�����s6��}�U�,�[����*dͰ��,*C:�m[� ��0����[9j�V��3�sng�{��!~�Fμ�_\�s���`��L�1�ڮ5k�R�<荔@+��"q�A��:�ꉿ�sm[��좔a�i]��[j,�q_l��$j��l�d�)E��J���ˮu�M���U���E5�ǂ��<�рt��QkI�`cr�1
z��<疳� ��1x.��F~�6{���N!���𬿣��U��1'g�cp���cCU2i���� ���~�������0)�jˑ��h�_���s���L�6�4�<��V�-�rKr(VA�Á/%]�B&�K
C��Ʋ<��(g�&��=�F����#ku]|S�V�|	�����6�1���0�L6��a{������{"�j�[>�<N<�Y^Jrvp>����.[����4�9��w-��������E��Qj������?CBh���0Z)�4��I�R2�"��;"�}\�3���5ȡ��E	��{�=9U���?`g�m
�h����CD� ��2e��ט��Um 8���c��Apq�W���s.#5�#Hk���%�t�� ���n��e����t��
��b��&����?[?�@Y������"Sc�6!_b�rV״2�n�YY��"s�'����9�&gg��{�ힷRfSv�2F��)t����O�E�D�\�յ��uUD1����l���rq��I�z�HsCԼ6m��T7D~Z[>���`���
�)�DJ�޺�>��Y�P�|I�.ZΗ�����$�=�πC-�L�+s��4Һ)��I�g(BE>NhW�����
���V�\���+FO�b�)_����7�0�KC�;�#&C��l�x�j(�`$�K�R��'����Toc��T!�Lҭ�n���)�����lbW�v+�ԡ6�������ѯ��0GP�B9ʔQ���ߋh����z����y���wM{b�rr�}�I�o�Km?IL��@�ܡ �uS0R֯�����P6\�k�Q�<|����/��v�m���7�*DZm.�A�ȉ4h��hm�o�SM�47���j��tr��
�ء��a��\�շj7��\�������^Z�wl�Ux��\i}n�js�C�Ǵ�Z_�	["~>��M�����5���,M�����L?�"Q6����D<�I������@q�1b��;��O�@� Yͥ$�[r;A�Mps�]ƀ�wN5TZ��~#ys�|X��cl�� +���	U�̼J�����o��"+�y ��8�%�.e��L�����u��-p�8_�ǞOng#O��NX��囍CG�W.���I�0�k�`�eU��p�U���&͇��j�dYǣ�+�Kp�&G?�̌[�΄��i;�`���.�U����Y���{Pq-�9��#�i��W�6FU���;��5s��tRˤ����+�l��>����q�,����sbX��1��~�;�����r+����!oc�*�Z�pLL@��Ẻ���c��p&.�`�q%@ʲ\�ʉP�IƐy9ty�S��3׫�"z�F+/\Yٽ��i�;�vu���&���цI��f�?�^�Z���/w��5 ��NɿY��_�s������ƾ�`��$��T^Ql�%Mh�taȈ� '6s{FcD|��i�G��!��*�S5���MDV�/��VM��.�d���H��O��=K;MP��b���eiӢ0T7�|P�٩ET���(�/�=���0���'��2X�¯)b�ԇW�k����B��Vz���`2}�����I��C� l�4��C��;��oB�)��s�?�lhP-��n�5N�z
]o~���zVf=���]����B�Z����`#�U���౮c�s7��~�|�2��!(O9K�4�j`��>����u�ҟ��b��,W�wL����nt����#��3p�n���`K� .Fџ �Q��3��c�5�-
U�O�!؏�R�����4�M>z���f��^cOq_1�6�P����[�劎x��ٌ�B����#h.0��_
j�?�z<�ø�rN:�ɾx��|a�z
���+�d�/'������e�bruմ�gք=��X��|ȩ).�M��n��ʝ����NYxp���1�\[� o'R|�A�|��8j�� ~� ���!�e�-e@y���S���i)&��B���3*��(��<~�f��G
�q(���Z���N���Q�� *�D�`�FQ*pҕ4/K��K�Eͬ�����2�^��H0LQ����vn�E�Y�X`�`�e[��".�2n���� L��kCl�au���'��4o
��wR�!���'��O���u+7�����y<������ķ�r!��fT�z����,���n����x���������ܰ���"E��>^��M��B���6�3��-�J2mV���4�'�hK߉�?*$j��M��<.&&+H��9�!yL��{����.V�V�m��7��ӡ7e�J�+��C�9R��(�����w�|�N���}^+y�����d��r������& �pea���Y�e�1h�!��n��kF:y����:��ĉx�H�P3��;�ֹ�}r�m럵T�����``l'��(��`�x5:��S8�����A6K!j���R��%�z9�D�ۇMAS9~���<�0�!���H=�e�X���)z_��0�ˡȟW�BȌ�)-����Wi 5�A�9�+K:�֖/N^��CBC�$��I�&�w f�0 Û�z)�كd�z�`h�>���{�F�)�qE��BRU�S1���#�a�1L�/=Λ[,�z�h`j��[$q�0gԀ���Ԣ�)4X�5RtǬ����a����ũ;z+��i�vH�4��8��iR�6��Ձ�b�nK��=�w�yQ@|Ć``c�#"@�T8y��l/�:Й�(#�Z���̶h���v��Aw������mn#�^��%�'R$Id�oS�h��VJ/��"���:P�>|��t������I�U��*=�SsO��Q!�1���.�T�l�(���#�" .����i8���ޖq[X��"��H�|��	 ����k�K��%c����a6&��D���.1)C�5���h����#|���9�}�X�r�)ͩ~��h�%���?��3�`�4����.�cF^��0,L���w��d�0z������8x�v;b$ʝ�:<��,L\q�Å����B�|*V�����9�-Z�2|��֏��~�H��
C�' ���t��p�VӉ����(��xsT4�Y7ʩ���k�E��j Z㋦���f��JyЯ��%Tv��5�������z �鎽7������]���ǝp��3r�  ܶ�4�d��-��m�N��%g�Js'0��$��M�uP̈���U?g�혗F�@?�ym��x�~��_���
��6�G�I@�J��X�ά�FK��
�r�h"�� P���."�)� ;�ZUUщ/8����7��>2�J�؆��CUAw�Q���"��w���'=sW�e��{cz�������6�ޱ8X
��X�{z&�'sٛJ��5�eOn�^*g��U��˙�)to��C_�;��}	+��M��� ��vi+ ��l��?"�+/���4�sN�t5V�|N�g�U�A�8�m���܆W 8˂�$06tӾX�W�S{��w�>�����u��R� Io�yhb����[q�FΎ'�y����m|������2��!�`8Ǚ�����j��^c��VWY�b8��kaѭ���Z�GO�<i�k�_p75��d�1�M��}5��?�!R�'��%�;糟�a���A��xYY�|���5iB-�׎���^��5��tT��?�W*|\���T�t�g����MHzs�Z�ʀ�˅�up׫Rɮ�&3u�	�f\)�;s�HC����p�/�G�A�p���c�ITQK�}���EfA�'r��H�Ҍ��&�2<�u�a6���zq-I�y����I0lEw����0�Z�1
"���Z�4�Jc�i�U���uK� U���m���\ԇ
��@O�
F�?ٔ@��TI3V�����8�()oǑf�5o�@S�eY�L^/н�5R�\0t���,�����k�E��^f�G Swa�2�^_�q�� ��A��H�Slc9ÚΏ4�7[��0�͏��t�;�zO�#[�{l�a9�`��>�E�$�f�4��9�`7L�i6{u�/���|����!�u���9�a,%^(oՉ�Μ�M����|n�q�`W�}y��	����)��|������*I�XЃ�hqB�ٵ�#�)� ��p�����4�z݈�A4@�d�nڗ����(I�w�qI+pzP�Ѷ����Ɩ9Rr�T8�㪻%��!i�RV�p0�	o.#�!G���1Ex�"�+m,��[�(O@���~6�z�J�:��G2oP���h��s�i���W(�u|tз�׆�`x{DIA�" R��~�F�6I��k��������*��jW��e(" IȬڡ���W�a�
݃����3ʒ�p$�K�w�:bV�Ĺ#�yK�ե�3~[U5�D̤� �JGu��(�ՉG�����0�k��No:!��<����+��U"�:}-�`Ⱥ5� bI��\���D�:U�=��Q���+Ez��(���+��RLgea	b�Mcb�L��]�$���T�CT%�k}���J[FƸR�7���=�gɺ,����qa'�S��4;t�SS�;H�;�J��=��#^vE��L�����jw�F���˷k�n��򪔡 ����_�ؤ`j{e�9�t�-fZN�|�_� ���kX��uܕ�}�6���`��X�op�Z��>��vaz����kr����#�#���,���`�%��,�D4ү��|�:����L�BǙnoz���=3�%V -K��hAܒkf�>`}s��U�||���|k��x̱�CkFG}��諨:�[�%���&�i�	� ���]�� ��j3H�H(R[��Gݙq!3��M4qMS��� ���Gھ�L��z�EA�%w�<�}����lӘh��S�.�dM�7�׀��ΎV
<������E2iLw���%�����&D��@���p�߈8}����C�O�	B�Uձ��5��p*�7�}����n��Y�7fQ�4�h~	�]��U��{���W�E�0�A�c86Ě�
���d\�÷g�T`�
0�sg��b��WB~�����g�~z�1K�%I��^]}��z@�������W��%M\��O6Sg��'(�5]_�<�Ζ`sn���T&Uߑ�ik�i�7��ܢ������ٞG�4�<���2����.;�p���'�+&z�@Rttl�})��B�tk F����y�MIt���?��?�@&����#�q����f鍊���6�>��`s�y*o�uF��G����sG�Y?%�NƄV���� ��渄�k�ng�E;�=���	i�k�S�K�4*�j����f��c"C�����ِ;��?�W�| ��/q�|��vQÆ��i�Sx����3:�l1-w��U��]+���9�Qy��'6�$�؁-_� k��`m*O]�_|>(�r��4AQ].�H��R�'�I4'���yS�����e�WjRO��9qX��lJ$%�
Q?dL�hC�Zn�Z�@����@ʭc�l����.�\����r�{��r8�a���6���)4��0�DxKؘK�|���gܽ:�>�l�����aY�G������W"����OgI�+�:�]�����T9�i&���Zf����qm�\#m����l��R!�򽬗ޛ��ˁ^}r� >4{ԍr�KYУ��N >�v @�x���d����^J���a����;[���	���!��!�jjy������e/Жꦬ�]�/~�XY���V����G�%�=�+'J��2�@Mz�P�I��������E�U�wA񙞅���0�%���~��8Ǩ�&�ZZ}_6�8�n0%��I����Ѹ��w��B�0�Z#�o�:la8j�ؚS~�� �]��@�En#M������)g+�IQ��<h���|���~ *�Y���V�L,�W�� ��@;�uQ�HQ��ho��T�]�� ����R���,ۆ�ee����Ѻ������E�����Ք��uq����b�޻�
E�t��_V惵��g�0}.x�n��d:7�(e<Slv����^�7�x�K��Ze@�}=�\9)kX���&bI�z���d��p�C`��.�>��S��u=�r�����kA/"��]�ߨ^��I�,C5m�$����7�ʒ'SD�*¯��t���x�R~nI8�~�N��:�1�_�c䚟���*H�8ܪ�|w�笖*�.��K�[�_�������5�9�tE*4$Y���F��ٚ
i2H��v�(�;7�'�m0�U.��s��%��%w���Q��Tk��Xt`�w��J[,��.��Yy�2���\ǒ�l	����K�y���;=v��u�@ّ٣7�g� ��a�;Ooi(��R��	G1?�������bL]��N����2�,/G̬N��a�C	�<�LJ*��;��� R��`�s�͹;NV2�~,���^2w� ޼�,�]&&W���_6�BIÿVJ��r����T��ċ_s��ǀm+X�:�	�)H�I�َ��v���L	U'�' #
�65��� �+�K.Y�챜yLl�
�,�"Tvυ�,a�.�Ȗ��Ѻ�)+C���'[�!��O��0�7�a`Mu�C]]l29���NTJ�WC[�×m����3�_��M�´�te[��'3��tKpa�eG�c����'؋�4�m�lQ�OxLi[F.Ên�}�x���}��S��semD�bz�WX*���s&�1�7�a�iLn�M�Dz?���.L�Zn�A����4RW9N����3�'O6ڠ����k�)�ֆ�����N�X؁�5{C`qd��ٛ�&~*���e�o:_:���T��7�4�����}��̑>fؠ��s4b떹/���^]Д0�R��s t�+ܲ��y�=	r�[���mZ����Y����b̋T~�Y�����A�La������J�vBSw�ȕ~t�|Sn(yp�]<j"�p5>mO���~w��\�ߢX�T������> yj�N�B�?(<�~��~�2�����pQ<I���ҢF"�hcS�'B�g���nj�UYh�n�rCU
���8��ѵ
����A"�$w���G��o��a�22+hJ[jo\����2�y��w{[o��V�g�B�rH���7 �J���y�::P��Ge�m\D�9��,��h��T���rpܞ��30��l��-�fۑaR���ب�ipF�M���"��4�Hz�<,��haX��)�ٜ���22����ܘ���C<ћ���F�h1��4L�R� �Up_6�r6�;٪=�f��?�b��D.s)�v�<�9c@�F���SI��qo���9�3^_·�17�zZw�p�dV7�_�J�׶��$����������oc��#צ�^$G�7��E�$r�[Eڊ���7;��� ��F����*i�T��"Qm�Q:��@2���|�⩕(��u�����K:��<U��L����@)���Gqϛj�L��K�,#Z0�-=�0R�Q^N�D#1��`�]Y/?2�����	�<�a+��L|�
����A�ν�40��.v< �����bS��Ͳ�-���vʌ�"�0�ȉ��pY~��D��p�{uj(ڌ�=�eͻ��Wu��4m,�S�-���}�����0��I���2�\�2~�N����r�(S��'.��rH�>�k=�ff�r/��
|Rk��5(���C3(�^���i�֓1�?�a�P^˒��,ē����P��.��)x�$�h���f9&+���C�����-�^�d�pr<��?8�6 �-��/5����v
��*��x�~�6�M�-����B���H�LA���D5���#�~_�ٵ��/�K�oݥD9u�����&X�G+k�o����JO����P�.��l�$# �������S�����fj����o�_��ާ3&�@�	A�?�^%3)�i�P�*���U3��[j�K��PZ��#o�jo�,g�."*�q����A662��6�{��q|�5�:#�zkJ54��K��u��]��+�r'��<��T'��^t�и�?�@�����%�����7qKQBE�u�(ԍ�܇x��;֫x��a��0cԘ`<�%P��N��B��R��I�&�
M��-�Q����=GS�P���iXO鮉�@�U���D�s߷��B�(�6���CB֗���2no����/����
��R�`�C9b��$j=�^�L�;��0��P��"�%oF��Ј�D�մ�Ŀ����SL�I�E����$J���%� p��[���K�Y�z�:�7A���V�����D��~����gM�4�<-��2<�x5#�Ǧ8m�AF�p���ĘVw&�?���1��Y��(�P(6����q�0Ē
Fg%:9�v0�(uf�i[ �yw��ä��í<��n�i	�K:�"�K@��UZ���o9�`Jd{�w\�Z��$���V�����1�*Z:�������*�]C�t�aد�'<�Ak����n$�B.�,od�R� Y�!�'�	W�E�
���!��
��f�ʙ�ɁC�G�m��d�Aeh{u�Š^��L�]t՞98.��z`%����5��YU(�%A�3*�'�W��+��"­\4�];1U� ������T/�&2�N0��\4��Z��� j.XT�Y<3Q]���ַ��"������l�s46�`}],�/��5	vR��:>,�˴*�xxp�f�س�,�IK�8�kb�`�l��:#u�p�X������;��ˣ"�҂����H���,sB����ֻٷ`8�_�[^k��+�q�F,ű�9h�S��r�A��mhX���W��P�?�zd�{Ri#��F���k=u���n�q��=�?�KH[B��vx�η9vu���GM�io~:�YhZ�-Y�!�R���������)�x��i���HS{Q0�j�WGX�]��nhX�~��0��3Q�b��{���� ��c�d��0gb�O �K��"љ���w�C:�x�I>��[��Z,�M��"@��O��eۤ�,p1�$E��^�`��fOgo�h�oɼ-���(�
�'� �ak� N��q����Œ��Մ�a1��+�l�]��5_Z������>�=�Q����K�otg����_]f�/�up��91�Ke{+#ܨL�1�U��S\�������m\��Ƹ��ݸ
"��E0|ERBW��0��-���[���	`��wQu��*������{S��¡��<�5����$eu[ �8!vq�Q��QN���^�_�`�]1]���H��C�l�����] 
���W֗#��P[p?{-�3�kD�AԞĥO8pn�2'�OUloJ�l�Jјȴf�E*WV���7V��^]>j�k�.�zԺ6w�A#��*>;( �J���f��YHvlM�����s����%|��5�tps֯T*�_=7E��z�g5�|��A:�� >.I$ثqWZ�����G�}����㒦����23�6������D���٬���;m��l�:	T�}�,�
���kq��1,Q�#U/o;ӫ"�籲� ���=�i7Ɣ6����}F_��1���F���y��\ ��"蹟��@�<�Ȍ7�������[��mç�I4���n_�oqD�z��;D64_M8���O��� �m�S Dn�M�6��.s^��k�����>׫n��G��l�C�$����ڙ����L�VhԻ��O�5u8��>�R� ����+����=	�M��CKH��P�75�x�2���u]�?�/�G�
/��u糏��b&�<W����M�mc�
mJ�\$"f]u�	`���� ^���X��(���6Rr���h�q9a�Һx�գ˵X�Aڕ���vY� A��)^a�?��:\x��g [X���処&��ot;������c.6,_��L3����R�:���78����T���|{f�0��9��z�gv|MJ��9������ZSq'��7�.�� /
wt��Rg��p-�\b�B�4/8�,�]O5D��m���a
�X�I3��2�1X�74�kџ�fp���i�8G��C2@��<�¤��u:��A��T';�C���,)M~io7"r򜙴��P�G@�XC/��.���rVsc�j�;U�/	o�rZI�?�4{�T����!e�]�����u��'�Eh��\h"���Z�3�<����d������9��ݴ���r1�5�igB���]��Ҍ����������M��������
j��&�EJ�E�Oa�s� �q�>�l�L0,.��O\�Av+�x(h���CB���P�/Y�R�l�+4�D��P�O*=e}a�����z�!j���(� p��8���)��v�.v���_%�L���A����4�Q�45)��˲�w�-z���C��cK[� ��B���R�ѻ$Z7����1Z��vZ����3^���Y����Խ{�O���B���n���Uٶ
��t�twѧ�m8�9������A�ֱB�}���e��e�f<�n�.��B1�5r��:O���s�ehᡓzD�}�:��E�\�Ϥ�^�9q����@}�c�r$x�,�d��_�7�{B��NI���b�o��W���jE�~���H�n��#�8�������{�p7�!6�]%54�*u+6���f&�)X(I7X9��J��ꜜ�;�_�}��Eo}EV�C*����`��_ꉺ�D�����S���21�<��������������f
D"48[j�nꏐV���O�n�����t��X}�ߛ��{��uy�����}�r�<'���3������>|h����t-8>
I���''N�z*�ͼґ;x��j1>-�k�����`�'#Moi����:�0�ي(}�b�FüP�s&�b-��|,�4��s41�c��<S�T�ԝ�
Xo�7�c�H�%/GJ��Y��N�`I���a'�\:���ˡ�xV��h;�${����R>~�>,��۾���l�)t��ӆ�$'5�Iߝ�z�o����1K���t#qm�����e7�xr���Q3�P��ȶ���H F4_UH$\ �Wq�Sb���V��>Ȑe*����lSن�Ѻb������{��ފ�`�f��p��AS,�؞<����f�@f��{3��8f�}ԕ����Oc��_ ���1e��L�t�
��0GQ��̕���f@��t�
B�ˡA�1
-������]��ܪ1چ��L�=�#MH]I���P����=��	��F�C�l]� p�˜R����Υ(���O6��l7����U ��Li�hV�vh�G2Ot���pY¥Z����i���I��z D~X`.p��Z���+�ݮ�U�:��*''[1�®{5���Pm�T��d%�j F�q��}\j���'�i�Pؚ��E���-�� ���U�u�z�~@ڵ��n��8����;���p�dR8j�h�Y׊�(�'K����[��T�i%SE�'��<L7�<� :ϥRbsϘ��6� ˡ��Z a�����^�j&�OYt��NO��h��������+���S�cK�'��~摍���vش5�Ԟ��S�C�|G�to4&�|)~��&�ۨ�`T�#����5Pü`7�C�˻�k[�I����4�B����*�+�����&��)�c;m�4�%7���J%=WE,`�#�Ĕ)>p��τ����}C\Z���l�����P�;o�?�K��#�I7�z��?zIx%¼vM~/�I�9i��O>R��h��w��M#�'+����Y��-�Lg����ēH���W�Lqc��1��P��Wjx���X�:`�Q�xݙhz��?HG<%B`�~��	��B��ыtP7���l0���ԡ��Q����%(z�Q�*e�m=��.������=bM��t�����Fs�>U���D�Ȅlj%+3�Q#X+vq���,����e�{Q"�ϸ�f���j��'�&��2	v�u�U�;��	ʁ��q��-�SlQ~Q��r����^l�,Aꔃ��n�iD'R�\��Z{�v�����t����к�;Wvʖ��K�����uϱ}��i��.��iw�y���(�&c�y��K�~c���|���ؽV��n�P�b�%X����|��C�=�IW��c�@�p�J2.�}!�Q����[i=���B�P�ǰ���,Y}��>���d1^�0*�7��	��-}v��%���|��/�y��+�t�uY����O(���_���7
�k%Q�s�Ҭcd�Qu�m$�e	�_�D���,:C�,a��bI@�� �~ׇP,$�׵"T����B��|�ө�&;D�x-]ruD���\�wd`%J��~i�f!&�?-� ��R�K]wi��+H� ���{�y�s�Fm�if^Q�.0�P�B$m��t^�'�+ ncV�YU �l���~�\u_.�e3���2\�maR���VnP���I��$6f�0�V��*���X��I Z"�
��/%O�e��c�ǋ)�{2�R�6��ő5��vP�7�uK�7���2��"��_x�+��k��V�\���u�Vؗ3-�Ig�p��}���T��UC�n���u�u�ݫ �F�����-S	��o���G�ER�Ӂj�&3����\2ԕB��lSt��2�2vG�re}��.*6��A;�TL�0�3�6;�[5���t�N�Bh���޿~�!O���.��!�j�l��������JwOU�\bG�	E_\�T -J�m�@��װ���ѡ�Y-FЅMָ_��7%���ܔ�}򬨠B��v0�P�H���g��l �ad���k"���%W�Ҧ{D8j!M���%BXF���~����*<�$O&� �GtE��P�0�X�����:�����D{��U}�Ϯ`左����f��j�uc�MK^殺���T;6Lg�>	������	F�F]@�[�L=���9g��(����e��K�}x�4c)]�Ώ�Qթ���9M��^\�V�2�}4�Y��?:���Njӕ����}#�� ��՗Ff��t�sr��_O��w*A_�l+4��A�c&���{����o������F�Y���a�~s��ȭh�h/��-�Q����n���Fi�qS�.�[?�Z�QS2$y���A���7�-���&_�f�ҟ"FaOgv�F��1G�8���5��o>�Eck��du�tT�`�M�hu���.g�wN{�c�������Ј� o0d�_i}��W���G�nT�SC�r�'�h�U"�g"X�c�æpK���ƛ�`��IĀU�)�V���?�H �:#!"F\!�j�^Pu�沓ƋGh����ی�l���k�Z���ۛ�������qe�����ΒF�
����/��[`�f�TI�y �4�t�=JoЅ3CA�	>���z@
�_��� �m7����C4a�c&Gx���&o3���I�Se�[a�~so)� Ea,N�;�g]��B(��>Z�<kF��5��r���Q�wh�l�b����uV�[;���ӱF�m�f���%�?�����p ��4�n\��<��j_|�1� Ol��֩��)g�>�m~���uj�Ԯ�(��I�Pp
�V����!ƮV"��|������XMJJ#X��hS�cH�i2�^;I6�U����Vh8�|2خ���}�hq=�9v-H���	Ƚ)�b	���o���(l�����r�S��J�YS�ģŴ�_�9���,�p(���e����b�*�z�K�����ĸ-8>�Oh�����ȩo��݉��"�i��$bʟ{
������(JC|�D�?Lz9g�m�Wݺ_�SY���m���U�c��nV��F�	��)߮�U��b3����[�4�0��"e��_�Pp7g�9Χ�?jG�ܓjR�пR�Xn�I]U7/��J��kq.{Ven�'�Mm`�d漛�	r�e/;I� %}aNJ�R�����L^rl	����ya�Z͘(�:�N�f���3G��d����Q=hl�8�@%i�sM�'�HZ�W�l���^1�Ǣd�
��o��B��m>�PT�g��C�3=4�W�����T�2���}��|8������;A{ZA�k���U-�b����{_����YD�>ۘ�hsLՁ�Jt����þ�c��jkI����p�4�@��\e���gg:�&���~�h�U����8ɦ�FUH{x��<9�A�g�����7k�N��՟	�|�ޖ
��N�b��T��l(�wҵ���N,'u��!�P�O2FXI��pf$t��!4u�G����2�d���I<�ψ1������QKkq�.�րW�^�����������\��4_�8���0O,��#m��o����&��܂��W���KH�;k�dٰ�]h ���xh����o^�'��P�33D�v趦�X��K���3e9wv5c"jaB&O���4m.�ǆD8?�ٿ|��fa���0Q�3����-Z(��Rݐ�u�Z哐�9��l�����B�C�(Zd7�B'� �C�J'2"J�DΤ�-,�$�I�+��}w�0�\fz��L��'�jN���W�m׉٫q.3��W�W@�F���S�:�J}3��*�yQZ�-��Xvl��h��E�[�%]�HΪT{z`(���!=aH��5�據Y�5E��)Z,�t���{��]k�Hu�6����(��]�^����7i�ԚVE��g��fU����o�Ɗ)�m��/��!����s&�5wqQ�B4��7����ɹ"��Fل#0vxu���j�����cBK��,�H���ɯW��ܬM{ʬEk��b�ZX����k
�Y����һk�Z�<ڂ�{�%� .W���8�I�w>�54�:xVI%l��^g(�`����R�p:��v���;%�F�rL��j��qNE��F���SP
�tk���������AI4�s��u�]Ո�է��W��շv@�%��l�~�%ێ0L��|���)��6�;��^�L��[��|�v�������I8���������d�6��Nsl��bݿ�}�
�@�(�d�{6�2˰x|$��a�W�Xsv�E�ٺ�vsS7f�W�FӇ��}O$&�P����� �3��.���@���s��k��u(�fHĂ���/����Ox��i��4X6;�:2+J�F�AK��sʳ�e޴4F���`c�1:pV1KO��U҅&RV.,��2�B�
�����i�KONR�� ɐA��x�8F	����r��ǳF��]>b�Õ�r�	3��!á�d��.��=�;��3eB�^C�d�?3VI!o�$��+����3����	��Bt�׳����.X�{�7j����᥯�V�dV�'�0fi�W��q;��AvNaZݜ��O��PR[�}'Y��T�64/"�Vwx�ʕ��bp�&�V�d\K�u/?<���8E��1���*����Ԇ��lX����v���j�Bzێ�:c��>,�$E�������HH�ʰ����X���&T���V��L��U��S��6#�\>��?)�f��FHa�a��)um���T�a�DEc���vֺ��dD ��#�:�z�D�ćOĴ�n�2js}j�p;��>�U3#=lt���"Oi��05͌N����`�C�U��7b��F�9�
T1��m�m'��R�px{OgaA&4�IM�9Ġ�c	2Tt[���\8_۱��AB,K��B��NMZ�u����ƞd -�Z���S%����6%^׷1"2���s9�޷��sZ���� �����0����Y�Ϡ�����w����!�yq*~Y���-b>[����N���iw�L5� �*P:M�ˇ&���sl���_�����i�(�;���o%*w�h0#��Þ�	�ٺ�P�����,�ƾ����(^s�[����J���&#;K�x�q®�.2K@m]���B>�'�i����$�p�o��}�n���ݻ:!u��9��ep����v,,~��ۿڬ�r��,��˺���Ѳ��1��v
���<��X�����:;<��V��Р��O�e�r��~�����o�)mV���:�RU�@ј�3��~uj�E��T�5Qk�����9�Z~� s��`Z	<� c�QoE%�-���?	xҹ�t��2+o/�A�K�<Qy���Y�Fc��D�<���3̲0�0���`{�*�TS��z��w��_��<:�����c�܃2˗�t�Rp�#���E���d�"�����T	_5X12+�gvz�ݭ[N�wk���**�-Q�
E����u*+$9>.�����)b�6�X��R6�Ѻȳˆg^PuĔU���J���>OM����&f#��L&���Q�ki�.ȵ��n���F�T�{ زZk�v�Nc����=�����M$a9�7���f\�J�E����}����_[�H���ǻ?��_�,-��9A��\�X������4�J�-[���U˹�0��M�육[&�OӚN���)	/
�s�(�O�y\$j���*�H������>�~"���r1��JK�c/�(s`T!8��y��?`�&��fVd�]^:�ހ���\�7�"=��k�JY���4KY���,K{�_��JLZ��@5u�K��F�1T�Z*��8���H��H�N�s���D=�����(�����zj
f�� 	"�y�-������T�K�֯�^ �8��,_hT����܀U�_II�Ra]�QЙ7+Ǩ�q;.d���:�B��$���\@�9'��@�{j7@�o��7e.�`).���=��F��x�)~���b�:�Lڈ]��S��#麾t{o��ǂB�(;^�3��]j9�r:����|M�K]_:f�Z�a���¡���{3��Ճ}X�
i	�����<�:޺^`x�'[l�TҜ���Up�O��Xx;H�M2UW�XC�B@����E���(ڥ��T�+�	�����w"�G5�yF=�$w����ʼ?i%[Љ��#	=��5�w�_bJA�(mEVbո�؆[�_����>g�Hxe2|�/��B��:f8t��2A��/ ��?����%�߉qH_]�l�C���Ś�FIJ"n��e3�)-��:����^Nߎ�s�V�|}������^�9���5�3-�Y�O"�w���c������vyYD,��2&�]�vV�~@�<ڤ���_��Ѕ%�]2AG��&'o�*eX�E]�,��J?#�W���ھ�冴�/��(-|]�;Rp����wI\7+E�<8sp�e�?O:�4�!��E,���mC]p��|�1�������js,ȣ�%���uճ�8�����GM� ��{�5�Z���,M �������o!ۯVd�e�IE{*V��Q��Wi,M�\��;3���3�EI��sԂ+-�\V�����Ou�t��u���P�8����$]j��md��Z�\���:;�Nm'զ~#��*l�POtlG�Z!w�R�)cUz~���Sb��8ǂ �Y]�$ ?ģ<a����*�R�j���X ��� �z/W@Qy����,B�3��v�����.�r�]�¥�9��'�hF���Y��2�u'0z̒���A~�}��M~�S��D.�\�Ŗkp�p�x�EA"}QG��¢E.�>�S��Q����:���ӞǋW��[)f� �i��&�v�ʆR�U�K�l�7������2w-+�t���le�j6��	60f���������3�Q�*烶��J���)�0j�%�,U|�4� �^��Y:��I���QZ�y�\��$7x(���o�^�y�0@���dTXeյ� YYx����(�/�3�nr*�y``�I�6m���{ɭ�)�E�.��QiT>�E1�)AzŅ�<CN ��!*�6��`�ăG	rj���}�"u�ɊV�XL%�"����9뱮"zt�~�n�тM�*h��)��$�n[��4E���90�;8}d��QHևhnw�㪄�������}|Ư�a���e�RC�B.CmU��#]V\=������C�+�&f����:���'U�s2�PJ�a`�����A����߼|�@Ğ����`��_.��Bè	�M������\�o�for-�~ڭo��"�F+<�`�1@p�z��փ�@˓�%vG����wN���{�5�f,�ȁ��x�@�h��C),��˼��䖯^��4W}�g5C���b���&j������2Mic:�����H�@���������b�u0���t%<�������ܮ�-y��.?!7F��`3g7_b�U��hdZ�x4���D���w'���N�V�eI�����R������u��` ��l"���u�m�F:Ćy4E�x�U��S#K��'�-�Qo��_$�.��"q��x<&��5��:�����(k�I��'�b�>�@���񪵮� �b�BЊ��@�����#��q=d�N�����9�mM��`�.������e�ǿH�3,xy+}Ӻ��$NȞ�R��{q����%ꯇ�8UҴ1�<�P3�X��b�ԇ�l��p�3_ƹ��a�'q�і.� 3�#���M�=K��� dd�2�P��^���SA���Nsc
�=���� �F�pF;�wjt��ߺ�_��୓���Ek����};Mxٶ�dPH�I�ftH$��O�^�P9��!@�'j)N�|��q�iqj�1���	)}l�M���\�S{�J =`o�r�ܞ�T�UIK2l�+p�et�S`��?"��
��ʎ��S��͞�[�,�:?3͗KJ�P�q+�M^#=��'�d���&�Y3r�q���(\��qm��n}���\G<��AM6t��P׵�Z�����u�^�XO��,�v��)�s+��˪zs).��9��Ϲg�_���X�Z0H�7����y��0���X�+���-����>���=M������n���#W�%� 
��y��͊��=���LO�Zl�i���J\�)�	��^�
�q1)�����Q^wT�p���>X���5m�9���jg|���9���e;���7�gM�[OV���c�����m�i���1��랱]Y_z����%�j۝Ox�<w�/�V(�EQ<x߆R�����Q�i��f}|��OrGJ�/���>���t���j�ϯ�m&�M�T����2��%n�3����lu)�B0�?	Fw` H���0���+�ru�!�X[���r�o�c� �Y�ͭ�r7�0ʔaj�dk��i��hN��r����j�Ȗk�{��'ů�5P]]sLNSaW��`":�r�Q�Jx���I̅��|�8γ�� ��'U�G1�Y���r�*-�L{�ٍ��a�>����B	Ou��\�q��8�)�*�m���8&Xfz�@���kD	�"��3lߌc�~�UY�:�9�^ҭ�cv��j�fuBa���Wv$ߐ��Ҡ+4"R�=>��	�h^w��Ɲ��7�
�uf�/�CyK]ӂ���_lu/�9!<��YC:7!v�+-Aț����zk�7��\W�陃� W��N��4���<�w�������G)�^{e:����}��]�b�E�o�'mxu)�ŀ_�����0�A|�.m|<�`[;��CA�����U�/�����Ca��m��Vʾ�����L���)��W�$�a�,6x������]x���b���/�9�����&�2ƬO����u=ϕ2R�ۿ�1�B�LҖ��*X@���J�>XU3�G�Ι]d�C�V����&�� J�\���r#���u����&��)<K��#���kq��9�+�`����" ��o{g�r͡�;r���W�J�#(뺊���_����\��crE"yP�Vd�e��l*W�f	)=�P0{�D�Ϊvv+�5q��i� �Gw���qޯ��՚]�{+F)��Rw|l�͂���:/�(<}H�ʖ�i�O@K`��S7�T�s��`a�i�3�|��G�;�"�F²3{S��N����SH/�q��sk}c��։W&�v勩+@�rZ�^r�R��xDN-j���ߟ�r[ Tf%�3&�܈����ģ�Ֆ�$���޸9�²b�����R��|�gjz�)�)\�j�y	���q���
�l�m��o]5�jK�T�,�ѫ�F�����* �rH4�g�rLe����G�s�ٳ(@��bA~a�xxP���"Hn�c�xR��Q"�Q`�c��HL�7IUB�%F8�%��Ń�Umpj�'�CZ�
�xۜ���O��-�"���ɴ y4,V5���{(�4/���~�"#���
�. �����������X�~��p0�-�J�`.�W�˔��u	C_߳مY�[>���
Wfeb���-��TSӣ�XWk���ƳGT�w�?�2-���ZC��cc7c|TI�]3o��Ň!�V��v7���S�(k�z�l	�Nd֠p�ֽ<S�)v!���`a��7�#�U�Rǻ�nMW�F���D��n��t�G(<_-z�ʴ~ԕ�s[Tg$�U�D4���}О̀�v�1S�`&VC��G��g�g��4��D��a�ʙ  �����33
B�'�?����3d���zB�c}���P�F��j[��s����%�#J�߿0h1��5� �P�vN�E�/b���������(� ���FA9;�n��
���4hL�����7�%m�Vu�A���]`	��-P����
7��3��+<�'����&"�L�۽D�ٛw(8.�=���ש�A�zI9��L�}�ȳ)L?Z�_��ա�.Z�[��I���o<���=���5 �O��4T�q�1%����Z%�6Qg)9��x� f!\;ȹ��c%eB&��I��l�����	@�Q�t+,�8/u��U ӈ��/�c�B�, �/�@¤�aq]I����\�*Z���UK�3Tʵ�
Y�r���e����L���nx.�;\�	�7��y&����G�n��_ �����9��w���N\pǱ�� 82�.�ˈ��⻑�U�ߊ<C�Ah�#�`�n,�L��-a��C��b�*��-�f�a���������>��Q=a�l������,f�"B���U�}j�qe$�dL�!<��������a'����v����j8u��;~X9C/с�������,������x����
p ��!VB¸�����F�#���޿����;��&�(�\������-�p���Ξ�l��>����6��/{G���|�3�T�������ؐt��q`u�4�@9�~��xw�:���P{&�5��.�TI��s<���cT=��1׉�L������(DU�O�aT��[���
�D+{`S�K��6Eҍ?�'�a+ �!�-,T½������h}O���;�dȨz�R>�=4 .�����m`P��ׅ�G�͠���{���ͨF̑0ȵD�0�`+�@5�m��;|Ķf�����W?���軎�*q�=kq��Zϯ�f�!�m��S�9����-��Hd�\Gd�T�c/5��x�9Z��E�̧������� 迖ءb]~y$LEP9m�qN
�CV��!�R;Լ�I�5�z�_��L>c�/�0M.�(���r�C�[[�k�G���
�M疼�<���
���C�N�`�W���i�]����u_�/�&?��|ag��S�o�� ;�Է����`��6(��8��S���S����x�8GF�p�J}�Z��`֥-������g�V���a�T�j��Wn�R��X~qq	��5�nd�r�ZM��Y�	K�'�w�v`��Y*�iM.���`��򣺮`6�
=�j��I�E����'��cќ{j��G��K��FE�p�J�5y3������ug<D/1����քp�Ƴ�%|�z���-��l G�ϥ��d��{N9g f^ܥ3�p/���n:�c54J��£�p~��Kӊ+A�)�Z,Nw)����<��� {�RE�E{�����&��zV�̍�*��z����sc����ŗ�s-!+"�'�����&�"��;���5m�v�̷�~�oTQRK�[<OGx^�? F@�� �h��������xt�/�����v����{����T���>�g���"(Yݢ�jT��\�e;`�y�e^�p�@���W�L��[�H�h3疄�s?'�	�:�����t@׮��@./P8/�2��d�[���w�;G�D��|>���3�=I+�����8j�W��KJ�`?"�?�a�6?�`��}�W��J~0Xh�b�-��P�$��II���s����
��@��w:%q]����B���� �2.��W "Kh%Δ~�[8<��hq9��y:4X/y����ax�����q��`��ϱ	K>�?~}3���ّ��Nމ��e-�P�]>|2 Nݭ&@�9�{ϩ�#��qU�׀�;�y�vU}�D��N7��d�	�"��MX��ԙ>'����n�=k�(�~c�;��q�d�t�0��ذ������8R�[������<�6tU�DG�|�����g05[�����D7���������W�6<���Z���.��0��4���	�@���p��#�*.
��k�#�h?�Q��5g��Mb������Z���w�����G����U	���mt�YLBcR>E��X3�g�X��:�t$A��������(��!0RpR�)lJㆼ�n�W�����j��TÖ��rnw:�C��^��=@�|.�x��ƀ�%r�������E˜)JO��=���a+B�>t'��6���1g'@�ڒ� :GЋ��B��N/IGW�����
�ߑcl8`(��r�I�I�w4������"�9��R4�cD���èZ�D�c�� �&�������8?�|I3�5R��L���t� #�>>-�V᱓�ء~�k��n�Un?r�Ѻ`y�:�[9R���ܞ���w��Á�a�y���1�@�SD��?����~q��)2|L!��ڌA���rv��3�>�����y`��2d����+d"K� �x�aR��FBL<|�+޻�/,������WW%�+�7Lɏo_y0N�P:��r��������%/�Ϳ�e�?�g����^�j3Њj��45 n��&M��"!�>��_GWb��l����F��yn�
�MIY��E����(�pU�c
�eK&{�/?~�zd�����/�5�ϧ�]�4�i�,M��,�یu�,�T�)�C5��T���A�7�WnO�vC*3�i���+��5$a�/xh��~~V��J�_�_3@g��'�[��Ly�Ž�慑��BQm���@`�"�!z�M�1�l�2Jw�8�	�'.݉�������\l�I3ˮ�\�M��1z���[��Óz��x�����#H�ǞQ�Hh�+_���wmK%Y�a/����{������R�N��\���푀�	 �xL L�<9	b�	y�^/�ۖJkC��ď�ݺ��&[�`�h18�f�m�>�/�dӅ6�xPDL=7e�[�Q���ȃo8������+��eELU���砐��t�َ��mF���1�#�s����A̘t�v�48R�o��[�Ki��4��۰�N��4�#�i݆v��Y��ۚ�ZQӎKH��[mՊc�\je�'���QZ��/Y��V5�Y>7����n4P���5o�o}����]�қ�
5��,_f��s����v[l�S>���ĄLj�������3p�A�0���ɝ8,8sD,O�����U���K����,vŻ��yo��Y�EVŪ�q�<8�S?e���3��:�p��Xl��t�Sh:[�2yt%��r�����w1�W�<[}����±��بX�]V�Q�B)l�
����Y�����[~Kr����υE�����-�iO�>�8�&��
���OE�?<8Vb����)UgE���k�M �>uܘ�'�e>!Qr��l!l\ǵ+c�t��0��N�Zs�]����uW���*3��4�1[�[�-=�5yo��+����v��UZ4��f���6�E���D��k�SB/"O�*p6AO�z�+ u3�Ҷ_��!ě���:�m�9"œ��0�.%�1�}Шp���I��3�kMM�[�/C�+�Z�MM#Qu���I��EE/���I���%�A"���e�{�$V�w��+�IgCO]uV1�Y�����*H�?(!
YD�|��La����B�M�v5�9~poј�m��T#�/V��{%`�5����n����/)�f6Y6{���9��#U��n���F�q�u��<..pp�-�LEx�Vs���P!
��^��̷s2�����D���v�v��bq���"B��iLP��J�	�O?U��Y��tta=^��|���{ͱW`��"�Z�ƌܵ��I%ar�Q����RS)T�E���?iT2���vX��#�wF�K"�q�\�$�ė&ڪc���A���K6�&��'�%a^.ǟ0��vuq��	���l�����^[)�2�+�D��F���u�f��_�����$:J�v�[��{A|�W�#�<+��~_'��g�E���xp��x���mV�1g$H�0I��\~�Ț^a�u�A��HBw�g#�!Jn��p�Mϼ�z�0��
-T�P�}�X�6��Қ��H�?�HP�~W�;�M�`������_��T��)m;����X�=q�\�1�ơ0��bF�m!ͷ�v/�@�j���&�@�!��p��љ�Ë't�u뾣w��M=��l�X�zX	nU$��J�z��{��ʁ�������97;1	d~�$���@�":; �����`8��� �|m�XQ�b�<"r�2�����%�/�I��
�q�4� ȭ��*�B�2�=r�� ��)/C�`tb 햷3�ϗ5=��q�g�����4�x��;���$�M��%�:����b{����	��GX�錊���������οX"�3�!8��f�)����������[���H���^����C3*Bk� �+ŤuS�N�<�µ��k&�bV�2�4̘���G=�l�Q�Y��ث2A,��|��N���ڼKҹ� ��):�zZ:�
�W��kc�(8���}nґ��g�@�J�Pq�Se�����zp��V���/��l��a����Jf��q���裉�[�i�kK%}Rj�R֨.��X��=���Nͪ<-���n��w*|��3D�י�w�*-���e��O��>׌d�e���T�V.�i��n�|���z��Y�Dj�y~��:��.�k��(c��p�@��!ʓ,ԣy
U 6�ۣ�l_6�������]�J\���6١)`�_��N*)��Oޚƛ��vהӨ�Q��|��!�po�=�Ӂ��i��&2����U{*V8�dpQ
a�����1��6�t��(}q�Vf:ua�<c���H�P���H�µ�瓹��C6��l�V���gi�w	���-��Y��Ժh�<�5:�#��ٻF��L�z�-:ÿ����K����n��`�GT�*��Vb8��M���ݨ���}ͽz���03�/9���n~y/^���U>S��X����pf�$t�a�t+s�*)>���*�]�T����^v_�L����/�	������䆥u�<��س�8����$<�C�m���"N��Ӂ�c����+T�=��`��@$�����܂(��M'����eXfyIO/v�2'�/y�;k��ꔊF�F�_�x���+^���l	_avA+I	��CFA4�m�'̿�ڢM�>2g�� ��b��5G@�)�C�.T2��GpT��C�r��0k�7��X;Y��C�`�j�M���@be5 5�M��)Ra_'{�����̵�㏙)��j�n�̶ rQ�RX<�?yB���l=X���v��ə����3��)_�_��u��g<���J<l:AG<c��3�����PK�/��rj+I��m�&ğO�����W�W���"��Hôy�[Ϝ���R�����/N����㧳�q@}Vd��.����c[����H�F.	f��kV���f]����P8n�\
��E���p�s;H��m-������$t���=0�ֽ�=JSL{�����]�`v~���&T:뾗B��2Y�s��6�ǁdIy�ZP�u�u�*�VŲ���O�>C=�-=5��?O噚�?��_���wep�ˈPφ��[��^��/��s����6��[`��gw�skt����m0սp�/#�F�`'�m�7��2(�BʽX�����ܠ��$'�'�B��Mq�T`G����p��J�(2���ܝ�y
8]~~�b4��(ɤǰ;�/[�s��Ā9���'eȇ�j�X�k���G��phJU�O}%u��]vK>�hg�o�\5�0aAu�4kx@y�jva���u���͖��5]��lAwm�.[l�w�QMP��0���)�:h���"�Wjiw��^R^���,Y�CD�T�!�'�n�����O�͡�c��5�)� Y���z����	8�NW�P��2��p�Aa<���VM�7~]��"ԥ8����Z���cŲ |�R65 ��f� ������>R��}�J�ۨ�����S���^�HC���L��^��U���KW�]�G
QӼ+u�z�|��L�z-%
�^5��.���BM��9�L�T�Z6�sӢxM�B*��m�22�-��[p�;��*��B�=E"-���pX�?�I2b_���ѐ�H��Ke5 ��Qg�����lI$>JK���/�`�� E�RحM9I!t��Jk�O�]�7�ܜ��j�Q���Q�:�:O�KVWL�Od�Q���.�k��������=;>X�QcD��~�ֲJ��@%"��>BQŔ2|9�ୱ�Ӷ�rR=l^����:ҮL7]�an�пX7������A��\�qJ�dUB�䈐��Y=�������8��@6���a�4g�~��6Q)��hP�g8m����0�i�;WC�M1�<`?��^����gDG�4���)4���Pf�(�A$�"9�?��'��?!��5�$O=C{nff�e-�6-��m#"���#��p��U1�'^�2�-|pD�d�T�2�m���zA��ɬV��2 +�A�=چ�CQ0��6*���]�
Y��`�"`ݾ�id�@�~q�Kl�h�b.��%	L�kF\�?��z� >�M�� S�͟E��
	��c:P����.Je�A:fO�;���aμ:2�S����)�GY�}��X�f�'h�_�|RdZ�����Nv��=.�1��t�eP\��+J�H�'	���<	�sȡ哊QK�f�Bֳ[�PY�T���JK�KE�?��iws`������Hl���ۥ��1�5Ҵ�P0�ݎm	c�='�Oc���< ��0�x?i3��8�W4B�j���	�nJiA���_ҳ�-G��e���G�Z���҉p_�%QH�p�/�e�go7������n�����G�_1I�͊��]���FR)��œ_�eN[-Ҩp���������=zEk���fw���%��a��6ϴ]ar� �r�t@�F	�x�[w-�)�C���
F"P�u?�k|��R%�E킦~7��N�;E��d�6��&U�S{/Q�	���U��L@)Ǧ�K�s!R�����\A܉�j)J,%�
�a��˂s^�h$0|�bԶ ��˂B��7�=_�+�v���Qﯤ�J -�;�Gs$C+ � �������0����br �����d����\4�%�zW[�B?j���~F͊ǻK`�fF�{R��qm��=����fq�S�%���hP���T�;�Ӻ��d}L$b��|�� 5����)D@�nV��n��>&�[�$�x���}	�x9����;�JZ*X������{���C�
"�Ȯ��gD=�U�bA��t��߄Kީ�j�-i�NbX孪~r��Ou��	�U�z���p�:����S�*?���0aK��J��J����������"�h��^m��epH�yN.:�{o��;$󳨒�^��_���x�:�y�K�iZ	�}�9���u��g�.9ը���,�E��	T��k�z�oO�,��_tb�}!m�����!>���L�P���޿�F�+�˚@���5~4A��L�}�[��'�%h�E��
0�>h.��'��E�g6 <J���h���̊�%��e�SsSO� E���Z�(x��`�x����X�H-�?e���(�[�����,�֐�o²��F�;�si�vo�zq�B)iמ>ONߧ�d�Ħ��d���y��?����h"�%چnz�|^�5�a���W���`/����L&��YCY9,~z��~��]q<�3;X[lJ�c&��U�s�
/�7�����M"$����/.Y�:`�O	;3�����5�������ݣ��}����Bj�,�#,�Mˏ+����q�"y'��S�7�<��ĸZ�ƄӼ���K=ϊ��J=S�|�d9,Ϭ:a��ype���z;q�$?7�"�f͇�h
�A:�K ⏵�6ke�ɩ-&�*h������薡�U3������Q�� �$�
*S\�v���X:sPlm����޻��𔲮b�$HQ���-��F��� �?CL�Q���U~�@�ީA����Nu�6�!�ľ>�Y��>P�m|�Et�E@�a�a�frr��9,�6g����B�|,d`��ո9�;����Ƈ�y\�.#��j�Z'�Tr�v1�`_�|��!o��)��Ys���h�Г����C�oA���̠�x��!x�b"#�,"O��@����"q�J��zpq��ٵl�`]�GUq��I�"�RƤ�̑4�������^�gY���u�� %�'8�9���5Ȅ�Z���R1�֠��~�W��eAf}���2��&����,x|��:G����i��	N���`��l<U㾹��.�ŝu�����A�/�o6����8h̄����S59'�ș�f�b��) z�f��3�x�e���N��c��E<���nS�É�r��XS�YU���-��F�CLi|��:àNw��G�
U?�s�/��m��hB�P�:�y�ǡ4�T�S�f�S��ӥ�f��z��3�PH�mr.�;���T���H-�xW�f�5����9�� ��=��1��c�{8��/=8����Ii˺��A����~�+Oݵ�N��Ў59��<3(t����������ؗ�:}"x�6�Gn��|��ɲ�'[���-i}E5�醪ؙ������m͐-��{��p�M�g�	k禍q����G��EJ�Ϣ�A/w��,<��_j2D��G�Qxc���E�䄶�� j�r���Z��PѪ�*
nN�T�Üpܗii�������=V��DQ�K3��
��2�~�j{�/�_j+w9����,�����!.KM�w�Ȭ�-��	�'��<�����1�6Q��S@����2��dV�B]I����Yʦ�������Ǝ�af�r叼ӄ����~�ao⣐�=:ۥ�I�y<}�����x$��4\ӑ5����$X>W�U�P��ߞ��壁���P�v����ª��o��b)v+d������CV,��dp�D�(�`�A�)]�<]��܀�\Ze�d�R�@��3�8g�o���tR����;͸�����L.e�����2ckY��T�;�ӌ���9��	X%h�.���i�AE��3��-srf�9�S8�9{�NQ�}�Neb�Ӱ��a�)�1��zЖWY"J<.�ܢ�
�5�^�~�ٰ�oW^Ǭ��e0������?������I G|�e���z[7��S��=�z_�77��d���^*�����/��^���e����BwqQC�1UĎ˶	_�9h ��p����`� � g�O��vM[s��j� K<�ZB^�h�R�,f�SqSޘ�*m�q�t�G�y�_�r,�/�蔞.�V��~֥�'T�
e�;�¢-�F@��n�)4�6lz���]�}�=ڔ����x��,�����h�j����s�* �vWN&f+�d��]�����/Y2�J�o�I�,��-����N�ׂe��\	�.�I��p| x�)�]�E�W�5��P�������f��P4��?�/9c�p�����yr�4m��$��|H�8<n���T����k o�
�ȝ�t������9��� ��jl1� ���V_Ό��|r(�jBM��]b���-��i4n�eJ���R��&5Ԇb
0�ˑ�U	SJ����S��9�	�����t����K@S!0ukl��V�3���m�C�Z���!Y�j-�	gĈ�:�s�e�o��6�<O�x��g����_D�-�k�!!R����嶄︾�������C}zM�Z	�O-&1��X��s �\�n�c�?]u���x��>�$"��N���K�v�Y�C����Շ�s&��.�D="3+���,�*�&m�0Y�f'�L�H���J�NJI��.�O<��I�sqeʮ̸VK��1c{`���P�K|���E�<�f1��_�$������<&�0�&^U�ܟ���� �Cv{����ư�ub��b�oA(�X}C�����]{*r-���x�tzZ�l���=�Y@��'�;roӱ��U���1_�)� �&���M/R��	'�Q��s"�.��;8�����w�R7����3VV�e�t�P�1��<#&��p��*�	��0��`M!�H�$�[8�_b}�T�Ŵ�W��Nɘ�&�[h��c�m�eش���zG*��3r*��>x�6I��E�{�׆��R�p|��$�}ԡ��S��-��Q����ݠ�8�h�Pe��m��3	/���@]����j��}uhn�iQ��2�vK��^��}W�#��6�U(�w�Ʒ0Y��^AΈ�/�E���iR(ĈNq��������gڣH��|���Jg�pe����B�aԤ8u6&��&H��񕝄._m�8-k5��`C�z�b�>��?��w�65.���@��%�5��֔7:���V���C�(3���8O���P�#H���L;�d��M�U��z1ȹj�G��Xض�� �
���Xw!�x�;7g�C�?���D�[����Q�e�8��c�	H���Wt�����"�,WL��dDϦn��^��;��M̴,�~4�L�Ƃ�itӿ���J�>S�Rg\�>�X��JJ��?�1.�+�LD���G��
qU"�ʍ��":�o��i/��yf�K��#TIY�u�VŦF��	:|���2�ɣ�oX$G�Kp��͡2���Ѷ���������*��ݕ��l�P
R꠱�c=n���I���ed����g�����T�5���"��y�����\u�D�*��r��ǂR\?puQm2�6����LV��A�X7K�C���QU�p���ċ
�[�.B�$�dU��~�;2z�9t�� �"�R�pF�E���^���X�\/��e5�瘝:�b�����^�d��C~ˆPbaZqJ�5Ѧ_DH���w�w�l�s��� ����l)"z�/���.�;�u�V��`��9���{���9����n�*��L�3�˃�	'ӏ���.�%/�q����"m�1�X_�cw�G�����|�#|�y�"��l�\[_ȱZUc��&�9?�E.�M���-��luP�Ĝe}�}ܜd
x3Ĭ�7X�D,^B��ڈ(Lu+ ���/+� x^�F�|�6�>��^;�lO)8
9�;�C~��۫4��6Ĳ�G|T� O���gK-��g,h6'�9�K���k��/� /�B�Q�]�qw��$+G����{4FƧhF6��7GNY�UT���X��� �">�ǃ�J��GMFHZs�ĵ\
���������v�a,���*��7��q���p�[⃨Ǹی��i����!n�� �($��J[Л���R��?��:Ѓ�������)�lAծ�Da^$�M�n�UXUϦ�Z�a�	�7�}%��T�f�ڲ�»���[
W7bʨݑK�2w���g���9Mx)̖��iKFL�ʹ�K���Zg	K'l�����-���AkJ�䜐�N�<��cz6h��(ߒ�}r�ͅM����x�N�X�fvj� �h�ntW�_�Ffk�I���zx�0�$�A�|&��]tc���ۖZ�4"^W�"���Ij�5�����Xd�e��.А� @0`z<�ީ�߇���A�b4�T��IQ{c�]O�\:6��`�����<f!����h�)S]Tw͓gf*�(`�5�(�;�&������Tpo�daB+
O�@��v�ZQ�J/[�	Vͨ�,�x<M8�^���!i�V��!O?|�����a��|^8 iG�-0����ҩ�2'?LyCa�;K�p���-��x�P?aD���vjw�=Nd�q�`s�����(nj �?�n�? (k�!9�\~����g/��7��g&�J�2��6e�R`��ʩ��
i�I�Nv���'D��E���j��L"���Ȁ�z�>�1
�k�e�XG1P⯧�G���䑌�0Jy���	� G��6�Mb�n�9VN�N4y>�W�8i��VhA��F�bV�f�Y��?���p�+a�-�y_�1!����@��%�O ����x)�[Q�2gT����E�,�(�z�L=�oG1ʇ���g=l�R:�	�@G�?<Q�~�f��#�e��'���^�V�x�L���Z���Q��Ȋ�_@1%6wЏ�'� �Ρ����9Ѡ���ȅA�fA�V���M*6� �I�/��|��
A�4����o/(�k{��*�--��복�BX�:�'SÚ&4�y7Ok�q�=�%�#K9�d��a��ą���C;a���n�8��i�"��C������\S�����s�gQ��.�bǸ�D�;S�K|��q���YQ�:Ɉ&��#��0p�Sܼ�
���Fu�@��k$�J찹֌�lY��)r��zT���'��?��"��"�<����j2#�e�a�d���-HUU����3!I�*���n�nQ@IS�M��ܩxƿ5٨�!��o�~��I�{�iТD����&̹��ݠa|�+U_w�?����xD� w�ك��G��@^�j�k�˨��]��c��W~+j�w'V��3�y���6v��*O��c��jV�±�d�F��]:n��k�l��T�č+R���)���������-/~�9lb!���3���b�)���j�c6�V
��|�s{��'�+���#�L�G��.������g�v����A�u����H��V�R+����rJ�K
k�=)K��t%*zAk�y_�z���:%��L�e�N��ƈ�g�+���qA��K��A�m,�U=�oDx�tHs����F�"�a=(���^��2��<ͯ�
J]�wƟ��h�#9��3���F��5R"�	|Au}@�.��`Z�:����>�_�6)�fk:r���:�
���ͨ
����h@�/�]f�DhכG�׳��a:�P�ZQ���yX*��߮un}T��;��DtL s��C��Ю ��n�[�\M��kSDTkh;4Ȩ�)Oow��xM����oϺ�	�M��HBb�A}�Ey����pEٞ"t�s%Q��5>I���\��=(�Rӂ��m�mv�W]A�i�c���{,��V��kn|��LaBFt�<S���xd���Nе�}��h�Q6����d�4C�^�6`*�Z�P0���Hf(a٤R�%�B4���͓s���Pz��
�
��H�6������/Ƞ4�}�VN�r`�E��r�TV��\�`�gsB����H�LB���A���h�5����TDN������g�	B�ܴ�z&貉&�L);@�f�5�IW�{�T�& S���IK����fǋ�ɿ �K�8, +r��4�]�5���-��P�� O��ch+�>ԓ�~tL����(�/=F�Z����7�o�=<��wH��\�!3/�n/�q�́`������Fb(b�a�ɟ��a�O�TE�)z*+�C�}�\�h�3^��5��Ks�N������۽����7�-d��}�~+}���$�܈���K�!��.?�PLI+�ڰ�Y��b+���i�,�tuj�JA�j��P�;���uyuH-T��[�1�&���m��n����!MK1}�L��.�`!�Qr��s�0����f�CZ�G�8��1r#Sx�?#Bz]U���i���2ˇ5��N�P�H���&L8����5�@��,��#l�&�	-t\�v4#��eRڛ�����y^���S��9���'��P8+W�]kxFA�Ҿ"�����X\DN�������#h-^�,�t�Q>l42*�YM��5�Ǝ.Jd�ޞjw�R�H�g/%s��X=�S}��]H�5�pu2̯����
�I+��g/��׶���R�����iǐl��BOF�h<��WQ�k$&zJ�	k�Oo�H��� ,ᅯveWF���'ϯ��_��+�s�s_�3)"|/���5�-]����m>�v�����֟+o	�������2L%��<���ڬ�!�{V�*@�J�=���%$�I�z� s�)�d4�w���V��LT��� ��!�l3?�z�YA�7�)���'�����;	����cҍЖW���Zl(5ȤK"@~Rcp�˩{"Ǻ7nȦ�z���cƑ.����C}�0L|�=�t���P��⼬����̊����t��6�Mt�MSԀT�e��1`i�'$��!d����A���W魫�<on�뗤�^�*1u��fhL��<!���o���5m��(�-i�e�@�O͊��f��<SQ� �E]� ��/�)������D���vh���3b�O�������d��I��֙��N_;��I�� ~濒67OY����V��uҲ9GQk*0�g	x���3�'�0C��	�깰|�S�2��j���J!̏��Ks,�;�]>��=�hτ�.H	�P�;]��j����$Dn�'D�;����*W����#l�C�(�Y껍����_�4���|H���1r�Ce��1�h�@��V�2���OH˱�{�Zų�{�[3�x��E@aUq�0P�{�.�H6�	ʐ� u��kl�ϾhX�:MOۀwe��A�+x�Β&�13�qM���U��@��m�[3N�"7�B+Ze������l��ⷲ����!����y��7ce�1�^l���������BƠAmw�!bjH�'6�b��/h�
�����Y_/jU�rSe�X��1Sx}�Ћ��Z��y܌tNI]* lQ��g�K��b��IU�j�i.cI���X��:x���qe�#�lN�~/9���/.qXf�q��%xuy�Um,$YA��v|]��f8AJ-�8�GrYg�,�����C�tC�(yH���-�v�d�u5�&��m�no�3)��Ah��OTI��v9(���8� 3(Y?�?�3�i"�f=x}�Š���k[Г���#�D�k8J ǯ!�w�ECԺ�@�"�X�@�e^�/�&������]���DpG��m.��^J����y�~/���)<>�� y��ǣ��]���l[����IK�������4��e!�J%_"�\3�4{�oރ@�W8�B(	��%�]2��5�Y3���n��7��k�5M�Y�|��1�em3�SQ�U������"��5�)�����Ը�iў�������,��Eov�AtBK�&�;���1�>�s/��4z���΁S���'&Vie߮2eG�	b̅�7�X\N�Bv6�9�I7�e�EǇ@!-ZX6*s��'.����`e}&�	1�I�1XH��U�L:H7�W���׸H�ĄωG���x�+�3Ǚ�|z�n.Gyg��꛵���BuFX䓋O�Η�1E��45�*���X�dŋI(C�?����H;q���.�`�;Ҧ�#h'���D#)��±��V>�h�lrp�i{����~��/�Mo�4g�'l�9^�����i��W!d[+��­�{���>�#�@�������o�	�gq������9�*���!U,d�6�����W�J��s��e�O�R ��y"��W����'7[xůV�A	ۖ�����~�-����\�/�u�<�{k�V�7�xC���Ӆ����$J�����s������3�]^҉A��E��=Y9��Ň�5�r�]�G�� �)�Y��^Ð�a2m�n̨�	�N͊B�\hMwщz���ooE<�'�f)�d�&S�`"�^]�Ķ���@����TɼNYMo����%�s���o�M�7�q)���Ԧ��D�)���S7�)��Qq��<�̓;Q�!g�;w`���Oz���Qk\x�6;T�r`x�1�ń��2�D��ZA>BG�I�m�k4���c��Ҋ`S�H�YRY+5|�gD(A���v�]�f��bk�ؿ��zF:פ*�Uv����M�Ϸ�B~i`a6���g�o�д ��4�
�^u�Й$�A��7��t�e��ơ����>R��g^]n��-�!ȫ��W�V �v������nڜ�>F1�E8��q��B��U;4��"��i��ׄ�gI�/����0� ��� ��X�~M��P}�	��܈��2I��Q�(E�:|`��>�9�,�XP����L���u���E�ϫpa� �R��|I�r7j�k�S��LHi�О��*J�H�5u�mh:CIDV3�����<�e��BV�ȣ��T�C�1z�b�-�I/O�a{��Z��� o,1������V�Į�;`�	�=������^��
Z���|I9��n��%��A��6Qs��!��fX`�A!�����9�&�xj�`���/��ڥ�$Ǚ�7�CS�&Y-�r��}}J��#�'��$z�J,��`,h>��K���b� ���lr�-�T�<�!7�'�0��5jQ�^��EF�5�|U7��hT%Z鰰Qg��KuI��=����ߘ6��J� XA@]�	���]������/P��x-z�q.�ـ�O)�f�%�T
��x�ا�+��7�q��K�<O$�2�&��Bp���zx�^c��+9'��]�B�P��/2:�T���ᶳM�2h>+��l�����pzخ=�D�Ҭ�
��X%0oNG��v!'���G[�;���a����j�)���6�6�f�a����DN8��S!@$5�+��X��5�fŁ��EQ)�w2q�]����I��*�L�sW`dA�\�U�$���:��&�	��P�����Џ
N�8N�B�gJ��e-ôb���қ�!A��9d��e�{跀�?Q�`X`�����(���^�*m��PV\�VE��|�6L�$0�u�L�%�H�����A�
̅G�:L'������ܸ^��56U��Qo�������j�{6D��ϵ�-9d��"ѬJs(�����ӛ���V��YC�`�h�1�O� rDK׼5�>������-��������A[�0�$zջ^�:�N���b-!�/��3'�"-�%��=�9�c���a����*H�r�є�0�����7�|7x�;�+Y�Ҫ{Aƛ�XK�.�	3���,��
8J�?Y�����Y�Xqou�dҧ�e��R���vS��7�����70r�n��-��]�E`�u����Va��#�R}<��(��s�.e��q�?D��Q�Xt�w��	C}�y�j&-�Eu�Q{�J/�iܵ�r?�b�(nzA��B
j\*��dGu��7�0�k����g�ւ�mu�'ʫC5��7��ؕ�6�O���eGhJ���t!$����G���ɉv�ؽ��W4�6v���Cp�oi����X�y���IW�ƨ&�IX�Nѱ���른�k,��":�h?ʗmxrP�x��8?���@1���(��)`��{փzŴ�0�e��c{��^c!i3L�֓��6�]��~:c��7~<F5�A�XI@g�;՟/��8	�x%�˕�E%��G�&�������&�|D=�Iu:6�$2j����ۏ��v���;��Z�1��D*�b6���9��p�����31i�=�W���V%� ��=�\��1.�$I�3�~���7Yi���s��³��2aq����sq&0O��6�Hb�H��q{#��3�n��Y������w=Ɖ����j6AS�t�����Q����@Z�N�����o,�n�ա����c=%�;m�@YWуj�8d ��/d̮�Vጎ���
p+O�|O' ��T���D�QkID���0�<ܜ�XK�bA�uN����%���5����@�ջ�X�-!�I�?4h� O
��f7��r}+V��s�`��^���p Gi������3�^4%V3!��Ɍ��-��4�M5:��?+�X8R�������FU��]�L�|�a4�/fb%�V����wڋ��%L��&��@�����U�D�����m�o�Z!ћ���ԟ/����*��!V�=�C��ӟ=H�!�8����>ߢ;�A����jK
_���8bJ.6?^~F�6��x>~C롶%_l.�0�:>�(�C�gh*ObC��)翂�L;~PHyB�����ڔ�V��%!��2_���
��fb!Ii@X�t;%�z�hs�����Wmڷr�.HM�}�)���ˮ}5uو'��	0�Ƣ���}�T��o�ה�XL���F�k�xP�>��p�ę�d�h����Ye�8d/7o��y���QR�C��k`S��Z�(m6��啤u���c�Z"�HY��jk���J�/�mZ�0}�R�蔊���~�m���)A�B!��-�_�'���-pvH��5��\�-ݦ?��g����A�Ɛ�i�d�c�6����� ��6����,�I�p�Q�Q8c�ּt�#k��-��,��0�@��@bh�U+�s�K�<��C��u#��['���W���	��z����O��M z��t�:4�s���}a&�J�.lu p
�����)j�c���⿭#uk;��,{����+3MV�U �+<sֻEC����\�m�y6"����y��!��hW�'-�q��`��f�޴M����Tč�R���?|d��G�2R�"p�����g!߶�PJ�V�(��yo}lb@v��=�T���5
9Cյˏ���߲@���Op+�0�6�/���q��CV�uA0VF�g$&��f�|�Ap�Sh��)�^S�%L?��J�t�^=x�<F=�Z��IvLo>�:SM;�[�)M�s8�n�fEa'vS���]���|R(y@^�jc��Lֺͽ�}�q�4���|N�O]����i�oG�3R�u0�ݕ{.��s�u�.���3����@�[3��ۖ��ܕ�]
�^=�2_z�vڐS8��yS΄k=�:o��Y-�G�x~��:��� >�eU���<t����Ľ�W^��RB`$�i��
;������ģ�rX�eyl�e����Ս3(��e�i#�����酓(��kcm�x�r{+UP��O�"ڽu��!t�F*e���?f"�O�Z���6<b��$ʂ�RsP��;
>]����S6Ț^Q ����[��fW�׎�/���]|~٫��?�Ȝ�������y��%�sB}u2}J:�+[�?1}�if���n�	��ǻ��u0'��{�>sH�q>.3qR��h���-�,#[��H��OXҖ�$��=t׶���Ʈl���܏L~E+�l�k�{���1 ��o�2}�J�H�/E���Sو,+��9Q��h���1�G�x�mPLI��ǝ�fl�",����b�jy�~7��Y��Ã��z/\z"��f̯v�lW�z��S����ڋ��h�L_��Fa�=�63n����ވr�Q�A1�a��뾜��F/�R)���'F����:����*2��4��O阌�l��ʗ���ق�����!v����H��"3�4E�.���7S��!�xF�F�]�Q\�XД©@�M�Z,���t)�;L/��13��j�f̂(eDg�o��.�`����
�<a����秳5���"��JqL�z<�9Ε"����𾄊3{���43�j+�A��:}7TS�Q����:�t#Zy6UY�������C��V�xT5)j�K��m�WóaW�����pSI�j^c��屔���[���˖2�%���wFuƚ�6�vf<H��TV� ���)'��a/���7m�"OAtpd�I���xE��؍=����S����74n}��F�`�б�^&c3�x�,m�R�7�h���D.ڐ�D�"�
x��~�o��K]a��%}�١�8>Y����>B���=��W�&�����c^
��
�d�&�%�6|�:ņ(�w��1���jS
��\=eխR���;Bn�;τ�Ƭ���i�	T���	�l��Ȃ)�h(u�.�M�{!�R"��lw<�p&/4Z�x��w!����p=������c��P]�bo�J<�ɿ�Py]�0B���EDk&Η'D����J.�"��4=�Ŋ��x��Kmoq���� S�%M{�[;J�Q[��*����/�B�P���h�(�[; �wՓ��_B �%h�;s��&}�SՕ���C�s�x��!b�^�p|jr���~>�^F�z��
"]��l`�y�z������J�����l
2-�:�c���$
]Њ��}��j�<�<���(�0F3��Zn����`n���"�"Icf�b�\��ߝ���h�oA4����$�*-l�[���;B=���h���N���q���v�Jv�3YB��*�����N�����w\H16����68b����[�sU=�E����V�4lZ�F{V�WaNt����Ը��:0�ɢ��)<�N�G����O~:�������J�� �Ji1�W��.��2��ps�.Z��tJ��׷|��$���c���й����8���)��Ӑ~�t(��^���<�Ki���I�l�&ڛ�%Hͨ�3���.4��>�sMQ�H����R7#���)Φ0�;�w]�Hi*
�fp.u1�X������qК��\�����.�3�2ؿ1����:�
��8�u�L�כ>#1�r������8Dh����,�`2-�5�G��o�;ʊ2{rӸ����?3t(���Ak}�I㛩)�?B����~�x�I�g2���>G���C�Q�&4O�A���u5�D Or	�]�G��߷�ޏku5Qi���[jmҮcu�Ʀ�z_�^���:�� <��k�BW���dh��IHTr����H/ۚD������:���3�if�fC��R�P���4Rz��|�����U��
�1�v�f���h���P���b$���	%jQ�
�?�С~�������ـQ��&��@�Q�%�E���,#�7�G,�����������tc1.�[����3���R��A�X�r�����f=�/=�eC���B�/�L��(+�_���5�JD�A�c���5�S���R���ҷ��^�K��\9k��%s� �$ /�������e{6ƺ���:��YX*,��C*��j-u@�xZ����R��+����X�3}$��%��V�1��s�d�Kb,�I�{z�T^$��>%�E�����̭��ߦ�s���1�e���r�+�Gp�ҁ�4'�ھ�Q�[����a�-aT��(w���$�-�Ng �S?@��b}!�6��4�ۛU�Y:j����c7�ip���l�,�z�?'f%.vX��)<$���o��P?Ht��r�:�����J� C��9M��Ѹ0"(|T	6�q'�򝮩��=�0�8��u�!ڋ�u��%!}H�e�fh�3u�{���Ol��S}�n��D.��� �����ִ9�GGB�c����a�O�m�W��*���q�3�=0o��_�E1�Yr����o��r�	v���RY��* �qz�8�X�3�2%����ˊ�s�=�S������g� �z���5%�+^��0kjԃ<;u3#=ֽ"X1�%�Yy�� �t�f�6�{k���.e=��K�m������؆4ǔ�v!���_�B0�~>��q���n���_٦��$��~UH�WX]�����pa�⚃�޷�ʾ�
��)z���bh�XD3ƚ�D���ρ�$���v�����N�u��pׯ���zW�o�KZb�R�˗Mi���Cs���u=���b�<��u�u��k1ϡ�=T�'3��;X�tD��̈��Lwhy���kнӦ�>��*�t�~�;�q.��1����rj�tԓ���qk ĺx(��L9pA��b�H�E��*k���խ<Z7��ų�fz��<�8�Ӯ�|�-����M��G��Yu�6�9����"hH�z`/�"O*I�i<~�Hs��/-`����!3a֊�8�b���|�	�ܕt�Lyfp���}�v������K/��B^���H��?~J�?Cŝ��E���Wg=PZ�?B㓉�HeZ2����3����v��\�uv_	����X)�).���{yD\i�ΌP��&m'G�i�NI���Zմ��H/z��?�cۤ��,��EU�!�����d�>�	VaE����Ɩ�
c�G��Ԯ>c
E� p!Sw��h�5��3?���w~���"k�,B�M�`�I7o�g�i�G�ׁ\�!Ѝ@ͽЋYF�8hg���A�{�Wް�x�[�=�t���8k���-e<}A��=q��5��f[9����#�7Jؒe2�s�~�j{�'[o��Rθ�OLC8���1��z	�f�ؑE&����A�|�|~>y%���5��0�L;vy2s"ՠ)��q���a�<zq�h>m?@��3+��"���<	*=;�0Nq����+m�}�d���X��4����[��%���!U����m$$��˿ڨl���(27(2�ע�ۆ���e�N�Ζ+��������Sby�tE7�	Z���D�.s��$X#�ѽcSLh$��m���|�e�ɻs4�>U�)����	4�����pK�
9fm�M���Tz:tZ�?<+�l :�)F��6�𰙖���$
�{��1���q5(��q��4�4��5f�2��F��o��u�s�`7��U�VS�rX���1���_�IC"�S���&�n�b��4l�h�>O>5FD8�5�P� x�*����~MR ��[¦�H�P�S��g �'-CD춧8�&׮i8(R�b�GFZU�t8t�.�P�pLy�k,��WǙ�z�zd M�<4Oh��/���LJ�2�E�daXJ-����K�'��5m3��
7�nǛiTB�)lr�Җc�����>t!+b)�6 ��K��y��R>F�C�N�A������=��f��z!Jŗ������,Wy�D���9'�ȴ�ζ�͕��Nи5$��u"w�ꪀ��1&a/�}B�~:��/!�0~{B7�l�d͝[�y#wU�^|���?�Ǖ�:�}�-�\2Y�0�Ѻ�3-�..s�4�`X���2)@���ț��<a�����m��D�Q�ABҝ�㪩�w�c_��|�� lr�6Œn~9���&�2+���x�g�d<�?������!�`�B�x&h߮����>��=п�p�A��@���AU6��8�#�դ�\��y��=.a�O�Xe�_^5�ݬɠj�fԧu�朎������^��i��%�f��g�UPkF���ng,Z������N��̨��,��o��|r��xSE��͡��hu��2Z5h�}�׍l�'�.�5"5a����O	���cn��H�@��^7B!儴%���~B����G���8���)qg>�WW�����de�h��o��p�eq�mhd��Y��*��4��,}�,��V?�9XT���13�D���F�e����S�����JD�wPG����W,QbH~��x�7��4B�F*EbS�D��f�Қj��D�zM�H��)�4�K>�Q�\���/nT/��\(�F�BJ�˨O�χi'o<���i�.8�H�� ��
���.
z	� I{Ѫ*}�%9�(����~���N�bZnJ/鐽�2�v̕�/P����l���\ؑX�O͎�lWOE�!K���Ĉ���©��V2�R>8�P4�ng���=�պ7�<rH�4���q����,m���8O�F��/#�xiݲ�#ϙbh�)TťC�e��ۗ	�։Y��˪�A�f�h��#4Q��Сx�N���n���{	&m/�*��G�b_��h�'�7�ۊ$H�ޒ�S�Ư���*i��t����J�[�nY�tpϥ��{g8}�3�>iiMl��Z�[����j������A,ݐt�c2c��7J�|�c�s�g�f�h�n��-5��pq�kS��&9�2���]���@�2o��b�cz��R�,Ez�E�LP89cN���xiD�1*�[�!��S���6���뗪L���������_���`W���r{V]�w3E��ܸ�D���_+��ɐo�׮d��%i��]k�:b�1˂��U���kE�ٳ�K53��u�]�r�'�J�K��|g1K���]��P�wڄR��Eo�ݙ�QX�4}/)�mr�a�� ̔��Uc�	���7$բ7�4^��V��5nd��
�5� S7��+1hW������*��x%asɦ�t)D#Y���Dͩ1R�Ӹ�w8w�K~��l=	���z���U�O e�b"i-ߡ��y�j��/���ZIQ,��H>�G�j�ި���Q���*�ezI.��D��yg
�{V��Y���5z��15p���:�$��[{@uA0��j�<��D+ A:c�!�TQO̺���Y�>nšCu[=V�_?�����o���۫)v}�#�Ե�{愍�ax���2����J�8F�k�(H��#�_8��.�n��>�1�)��k(��������Bkk�x�	U�(��FFmIH��I��!�*�Km�`�-�s��'Q+q�	"��{��{k�C&h%ZaB0�~:,:�K�x��H�1i6�?,P>�Q�!�q����]F�r(��.��s�P!��|���X�P�>�s�gc3������=��2ޙ�i�H���C	)o�X��f^�r�uwB��Ť;02]R<
=�_%�
����̐�#9�MoS�S~���qe���w���/P��-�Y2���?O�������h|W^���m(�$G�1oC9?0�#�-_�f���n'�FV觹o۳	�6cV��8i�d���t�d��B/Zg��KT�&�bo>Ҫ���$8�3K��Cu��G����߾�L�͔  �4�%9�>�������F�-D~y�6]c���=��'�A��B�/J �+Gs����E��Ի����.�ڰU��ޟpj����h�8�Q̎u�*���<�h���3���f0�P>c��-W�6�y�����Ѵ��b�'}���5�����*0���fl�(��1��y����HK�6��X�)X~�7s/��!���nyV��m�J�_���Ie�iu�ў:E���;��/����x;Y�&��8I��D�;����ʙ__!�e�bu��*&��Ӿ6�������V��s�Q
BGQ����*ě��WUP��K��x��������}��m�ޮS��΅STA������������\TIK��E7��TJ���rJ'y��vp���7y��A8]�f�7�2J���A@����� �)C�~v4���d�|"y�S�?o]�=�2�ٕZ�`�x��{|����,�u�)D��	���]�@p��b����B2k���̑��4%+9㘤@b4��f�!0:{����>Lf� >P�v7���N{5��H�M��x��u��_�\��	�,jL�j#o��Lm	N�.�$���Y-U�n��l�GحN�25�k�K"�{t����[���s�=�����"��|�h���r;��q��X%Ԯr�ػ(��5�Ƥg�!���
7z�o��'�ԍ�&Z7��3�C&&�Y9�4��=�R2��ַ��_���)��
,��f��9���V��/3��z�=ʐ�{q��.�艵͟���q�1�G`�غT	p�`����^|�~��2hZ�Fה�R�������� =�?j�>ki�`��*�	6�Bϯ��Z�`-�!��ݿ�����}�{Owj�i2I��ƽx�ķ���m�Hn~��Uٛ>�c�/� _��ZFaɑ���f��ǹ�@�Xr��)�B�c�'ْ�룻��v4j��JQ�AW nHtm��e}-@��o��Z�(�e<����z*�/.yp�������������SX0DgD�uI���|�1�i�=ş�� K�F7�F�c�G���ق�f3��D�zG%hyԼ>����`���(����ىs���~{�1F0r����kf�����4���_|n�=[S|���}�&{�w�xfU��m:�'%�r4�PxJQY�wzkýP.�s+doz=�I�91�n�#����t\�D���YRWå��V�3Jj_����W ��(���]�H��V��^���RiQ.�$����8{&&�şK׎���Z��K�Y�E��J�4�h�
�k-[� F�z�t`�KI�t{���Bm�*8��3 /<��D�^��U��rJK�7I���Vi�f��/��n�B	��Z�̳
��f���=�B�i�ɇ����+
"�y����-1�_>�MX����o��M�X��Bq_Ҿz8��Fק\_���8j���p:䴡\���vנ��.n����g��#�ox��4,�}�Ⓝ"�6�r�;�[��ߒ��F����ȄF��K�ԛ6�@�q3%#GK��%�"~�{���^;�����O����8�,[��}�x)��4��E��dg�y���[�H�3�����W԰�Xu[��`���/��V�#�pQa��Bs�04 �?MI@�1�ܔ3�s�3���e��Y�L��o�i����8���&|�H��f�zx#�����uy,M����8�P��r��$r
�e{}���s���N�@�j��b�$��8_���C�AXp�������;q�2��5������dE���Z�_h���UY��{:��8<�!0��iq
 ����S�����>Xg|����W��.�Q'���������j�^ZL՜W��U���h�8���a�,o��tgsh���ɺ%������q�p��V*��9��,��.��\-h�P���ey>b���{�]���ɉ��)��]\j��/ju-Zޮ���JƥM�HSD�v�>�O�%�g��&����ӣ�j\��Ɂa���*�5ŀ�0��	}cCi���^u��Nh�g:��c����w�"�m<xP�x$�\���(���b���A��BީA��F7Wb�X�� ̢yM2;gq�U��V��|26��k��5�k.J@҇����像#��D'3?pk��\���aC��ݽܐ����0/e�7ZF
��|��tzK�E ��ȿ�"��d��*�3*i���H�Ȩ�u<���jyǤ['=�SW/>MԨ},f/<)v�#x2�	��Z&Y�M����SG"��PS�[ �����Y,�0^/<;��'R��D��Q�3�z���i�3vbލ�����%X5;L&��n�ք��
u��� �7_YE����Έ0�T�@玷��	D$��z*+��n׳�K�|�]3�X�C�PR҃>���Ѩd.H?E�R�T���z�^S)�� or�U��w����S'�hj���&�Yʌd��1��g^�w��Cӗ�p�ąF��<��[��a��[ q�L�w��N��pc,�N�p���6�z�Xi[�ȹ�W�-�<��:�7
�u/u�A�۷����3a�:l���h����,��dN�6s�?u��3xp�!-�LLz�Ӷ�����g��<�����>��%D��������U0#�}���~�ݞ��ҴxO��&�!lP5(W'vt�$�r��a�����W�n����d��n���Ҵ��lF=8�%�%�����:b��l�x���
��o �ئd��'/JQ޶*����{A&���><AJOVG�`D��/��^#9�&ע�oobHh(�U�-�ԛ^3�����$���8):��E�Gӄ�����T4��O�׏suܑk��������cU��,�B�A����Y=�1�]�p��дxHcC� T����/�����η�[�kۀ��Fj���)��B﬿�܉���qr����gs�w�2��p��T��]o 5LvD�zCvK���go_R��x������|��l;���8���zj���'�?A?�b���*��O#�0�S-O[�����a�x�������e�-x��-m\�}ж���j�ۆ]]�)����3y�Th�&�(n��B�(("�v�pv�W�'GB1�\]����R�G��{��
��$��Ύv�룃4�ְh\�E�rq��++Z���u�ڃ�d\�KO�\pov��K]1��1��e���Y�b]�]%����uP���rL-`�K�n�|����y��s��JU3�u?5�8O��:ؔ=���2d�6�}�,�Q�-���7���c���~Q]�#�j0=_A�X S.�P�'\��~lǪ]�7 k-ЕR�L�$��W�����g��#5����K`�7ʮ���Z�j'��*�edy��\�K����������T1��!`n΍��xU�t�z�D]�
U�+q#,�O��>~,+��M�\�s���O�(O`�,�	-�<N��N�5��5�* �+�)���+�u�Q$*U��q��
Q�H�.�j�Zfv������֦%�a��� iE��m���ݟ�W��~�z�|��<����$4��_|���q�wG�
��^"<���U���9��~#���tX�/y����[�ڔc�����1�U���xÖwN��מJhU�'k��g���q�[u�"W���y]�%~)��˃x�`�lA�'癡�\mw��p-���JX� wH'��!
b<)�uN��d^���0L&|��µŰ�*O�"9M��t������4 ��Y�Rϟ_�-4�RB����c���	/m��Waϋ>��W�4��9�)N�1�:
��ZX��0�_�Iu�k�Z�(���S��S������[���Jc���]m8�J1)����D@����G�{��pG����5t�gf�NG(	�,����X��'�Ru���f���l�t*��aD�T����t�J=ᦖ%~y;�&�����zs��H�i��R":�������->���Bc�叉.r��3�t}�������⋜��r�Fe�6��}�"GQ��!r�e=�K�T%MÔp(�V�G��{1��S����j�'Sh�0�Y�����f�� ��I�k髀�2Q���{'��q��-����`�U�\6hUM6k������׿��ܩ��VM�������V�/��I�du@?O�e�"#��̍`>�k^������,�3�GW������o���ظB�]�vb	��A�	�\FPz�EB8�������]e�"W/P���L���og��Z̉�@d��a4uC'q��a�IIK�GH�:|