��/  �(e���&��)�t�����RĄ��Z�q�O�?[���ӓ�w:�~�*A�0#
��:o���꬏\��H���m��"��L����.ᓮ���B��W�W&{��Aa�(Q�V�9�Fo%׻7Td���� �7y��=P����?�����Y�e��,�	�^��<�J	9�yI۴�:Sހ?�!��mbH3.��^;�b1�A��Y��7x����i~?��@� g�3�__T�םܪ�"�|�
��bwO};��9���G��\�l^. ��hu��ny��~�2�`�/Q�z��r�3�:�S�[�މA^����. w>�^�N'���[�չGn���'NJ�H�7��\��|1�iįI!*mU7Jom]| ��W:m��-�j.T�g.���Ά�;��~�@QrXUBY�A�1}	�1�+��R�����I6M+*��� `�������҈����]K�<E�L<������!�e���H�����(��M��u��$�7��2wľ�UG� ��p�]ܵ�~��2,h���v���jE̶��ۣ����'��f�k�!xV���9�u�a��0���w��la��B�<�����"?R>��s�>m�ǳ=K��UѤ��y1�y���Z'��6l�����N	�L�i.ӟ]� r�M���^^�U�]"SkQ��(���㫵�p���ԔF��ч?L�]"�T!�RC~��s�!�L	���P*�z�-���KH8��6ɇ!��-f�� G���3����W]U�ǹ3���x�՚��|Q�)!��q]Ԑ���H$�-�/J��_ٗ�V�n�Z7+ZK;~ʦ��y��E����Ɠ.Yy3�L��G'e�o*��+SR��?_ch*k��v�����Y>R�2���!G�����5�������H˩�(�;u�X��/��yr�a��D(:xJ�GZjUk�iQ�c��^��A��v�Kѿip���l|�����PĠm��B��eU\ ����Y�v��kJꚇ����4��]
"�WE��n6\�"+�"ٱMp�O뮶��A@^��v�Z�h�)��]Mp�d�ĊÌ��~k'�KA�j����펔�������]��E��*�:�%7ò�l29��M)r=������&��ig�o�e^�B	���Ͻ�z�f{Cd��]�<ׯ$���&.f�X�J�p�k�f�NU|�D-���)t�<���)��v��@�rUrq�8�2���Yda�y�f�э��LR�����Cq��!�
�Gw����A[ c��ݹ�*(?���T��?r���7Lz��,�疡n�Km�>��@�h��U~$,6�s�i��[�EF���1iT�84M�5�5
��[(;��{��V4ĵ@�aM�FyKƖBJ�L�(��DJ�� y�!���ӡ8C3],lr�+��ɔR��l:̜,/�~J������m�����N�����"�l�' Q���.�l(�#9�>�ע�E�D]���.�]�c�_�\�gj��X#UqMA+>��L=(s�y��Kˮ��!��ڐ����@�]�LBm'�{���MȇH�ml 3	1Sv���5���%����kW~��P`��뿗���,j��������Rm�6�	��x��3�!��,��K����K�fs;�o��ϫ.��	[|���K���eK�	��O�":_�����0}<ɬ���w�.ƿ�O�W��!s+�c��+���L.�F�� y�"<�˭�X�ظ~�[t�6��AB�"��-''敀����_�tw��f���.�Z|?�����"��P����h�$;N�	��Y�?��Kv�
�GYW'��g�J;Z�a�;0*m��v:��9-r��g�*���Y��?E��I_�q��u'\LJ���?�r����B�Ŗn����
��g���Ç�yk���L3F��aD���i�v�2!�h���踮�7DP9���R+�Y�EY:��C�1Y���e�X���,:�|G��eW&�d�3�W{�����9�+o�\�QwA�����om�~�_��_�tms^��6��d'r���
ۤ���Ǫ��+���NN~������ 2�E �u��W�[�3�8�Ż��q."�ř��|�)�$�������
`2��:��j[��SQԍ��`"$�~��@=:�p]��^eK�^m����R����+�T\kɼeՇ���+m��n��dK\^	��t%��O��7�<���(zn��|3D�ad�A��`oZ>8"�A��U���"`��eu&=$ٻbѰ�=���h�b|�`��;�\��$�2%����ПV�Y��1uGPș������"�gMPJ�I�"{$����;��:72=����T�4e'�����R^E�P��n��9VLT̝�����^�����-�6&���VB\��ݜLS1ItF]w�a)lu�Yh�YQ*)��/�-{����ևpN��+6�s���ǾO4���"���n1QZ.]0sq���0]}M3# F�g�Us�8��.DnVK�����~�6sޫ-Rn���O��Swd롟�r�JC aa0���]�Mc䢃* `�Qp(��4�7WD;}��H�=BǨǐ����ˊ�.��*Ѹ]�6Á7�x]&vY�8��c��2#�ZO!m�B�6�q����N�.��U�����h����x\���Y�W�����H9 "�2 ����ܾ��8��t�\��oDO��a*y�>c��.�]E�d�y�Hhi����X�h�;���:<`A�$���^�o͂�Β��jl�}pn�]'�	:rꜥ�ZX���I6�8������u-����+$����8��>���<6ѐh$��N�U?|ޥjKu�G�/5O_��i���U!R/n�C�$)�L��a2�Eӈ@Q�Ư�ֈx�kcTi��#-�&Eu���g�"*�R�8�'_)�(
'�(��r�TD�ܛj-J�m�x'��_`��r�� �7�����IF�%�c>yǆf꧹��޷d�K�+cA0S�Xoz&�7��O�=l<��0dQ���n�b��g�c�qH
�D��AZR�#�U�)+$�������$D4oqtxq�j㔰òR��;%�.yl���"�!=��q�k"�a��Հ�tY_����ȹ����@����P��$W���X��J�N�z'��RV��|��k{�G�׀����AO�5: �g�=���������:�_���ȷn���0�6�RH�{QPM5��9r�S nƀ%��}$�#nS:�{�dr��Y[��%��)�@E���w�Z��c���̗�o��k阑⥻V��*N�� ��Fִ�:�+�Q�"aZ�7"������i�_�u��'�/���\�[� �z@������yO�T��u��;+u^�@p�e}�bL���&
����� �u��p*��u���LǦ����2m�:}��.�4���$��;�qU�^n5jӊ1~iX���h+U�-�6��G���QJ�>��i�~��Oj�7q�M��Gj5��cB��h%C�h_|Q�����eT�����c��N2C1梢uy��m/�J�S=r���ӕ�_1F�e��2>��{�M0�Ң���e��O%h�5���1�)7@su(����>��l��	���[��?!��TJ'J�I��M3_��fC9:�hvU� H�����h��C\���]ͦC�8���K5��U�d)�Q*"��@��Lt�0�|�5�*�Rs�9y���C~qBf	$aX��rc�u;���o�d�@�(�ow�#������d���=�(	љ暵�� �P,�@Zi6˯��r��%x�B�NWvT�o3VR/7�`c��!�^��S�絎85�r�ig*C�0H{:�WG\R��O��E��K
�pn���	/(��zkN�O��G�g��1�I&��~Â����;ւ���Oo#�*�Wgq����F���V,��{sj�T��U�ë)�\"�:�z~��1�ԃM�+����,9�V���x��s�T��դ�|N��G�*��"�Z�5XM�X��x*%�4Wq�
\V������/��e��%�^�޺��e_=���i�Wȉ��F2�,>���5��ՔF�)��=�ִ���2�p�ܐȯ}���v������;�%�;�a~�V���6��	��|����h9�vI��H�Vp"0����t�M?́˼�oCV���?r���l A��\�����V�s��k�]%�]�띇)�
-�Dk���<7���.�!�2]I ��S��.���L��q�U��*"$�d_}��a����Ă7<�nn쓠
��JOp�N��2��kv�� "�m������D�s�+�d
2@�B�Ud�����?(��D`5J�;;�E�?�;慦'jZ�K��`��G��-�f�*�7r3qf%Z& E\�c�Z��RQxB���?�]�X}܃����	޴�!R���h<�� ��S�&�Gz��0R��r\z�=(��	���=��es�┪_G�ρ��,��=��lg��1�}s�	E���O�~��&�W���2���"�O2K�ƅj������i($�y��aH��taM�<Ҳ��Wv����s~�
*z��K��b�
�������W��!߱��yWf,�2��4��0�V�;� >54?��.7�$\@�mʎ63'�b��y�st�/`��̘��E�������7�֢�1�.�Ѭ�֙�G?�v�Kv��8B��
�Bf���ɲ�c
بK��'P�����m��.W��<����L��;8j]�{�rŧ�N&�\���Q�i%<b����>E}�o��-C�g��i����Unq�Y�G�僳\E�я�p����zd�n�eb�.t�7��� ��9KsM�'��?�N���¦ᩴ���F��JX�,�����'��+�G?�hM@)�QH�=LC��T��Bѡ����cU;��m��@ͳd������_o���b��b�!���A]S��T��ʾ�B�>��N�Sz<��no��?+m���5@b��pyg�jQia�F�yڝK�z2k򀛜�=�fHXC_�o&L�8��no��EX��r��C$�6{�PE~U�T���"�z�fs4-�g �g͋70���{�ŃT�Y
u؎tGL�,�+��X�dשWW&v`�p*)}��C|��y��4}+P�SJ����"��oE��� �CjZ��euW����F����`��3��ty�o����_�&<�/Q8g���(�Le!-2�&2�lcZw}"h[qu��>��sn�'���*x���Yr��u�(Ps�p��������ncQ|Na� <(�tM�~!У�y�k��1?��Ph�BSmr���=����uݰ�����}��V����V�����U���Y4��ׁ��ߥf��;�:a@���"���l5���mî�(�W[�r�ا��5�+�߳�L����(���(�B��b?���
ey0"��u�:vYo>���t�����ͷtk��aJ�o�- ڀئ���t�p6����e��/��	]����U��:�`�w���@�ƁL[L��[�z��
�W�Ԛ�at�`c���P��N�"0$�A���t�R��~�T(�ҳ��'H�O"G˨��֋�q�^.A�" -����qJ���MOQ��R�b5��u^B��p'Gr��kt����T���yU�zT�\���׀'��[&Nͬ������yh5:�˕�]�d5�r�%?m/��%
%��(��>�V��4�֢��6���]�ռ�4�km�/[o�H@*�?Ӛ��!zC�p�}��V��y!��Bȿ���o'��y
a�iAXܩ��u��p�+���WJ� aŮ��+��Ӄ/�/�%ĩS����5��G�U\��52$����i]�tzYxD���4ɼ.�a%������H�R���m��%�Yx���N|3}���e�+),rL ,|����sf�Ǡäڗ"y�GF�'���di7Jf�R�����//�"�Y����C�&��c�lq�Fk�bV�y��&�ln��(��f"A�]9���릪.�3ԍC���n��t�!qU�S�V�"�P��$C��Įm�������v).'���܎�I�*S���]�E
z�l����A���@ԍ����'�K��n�+���@��؁��k�+?�A �d���L�Ux'F�0�L�;�X�M�.�%!�0z_�E��Cx�/�K��ʴ���ﲪ���7���ra�mg���D,D`B�4�On����Po&�{H7���9'�Z1����\�(�!�YCȒ���0�ғ��zǰcV[{�ҙ��
i��/l#�n�7�Z�����h�5a�w��ˋA�k�(χ�d���ʙ�l����q�,v|8�-ݏ�Z�/p�ia���u!K�c&C7�O�IvwG�a�sŤ��xy�@|�5f

w�n�.0hAĥ �G�d�MhϮ����G�د�9��Z����t�'Z��+�`���a��f��`�^ZPP��|�ME"lP����Ǐ�s�J��>��~)��W�՚$�v� ���&*�$���J���� r�q\F(���.<��	Gc鏶f��[D�������U҉�@���ø:s�&/3g��+��jXVMxr�VzRfo���[-,Q� ��#p���y��Ipx�r�[��f���qqӾC�7ܒ��uK����ӻ�}O�*9�g����#8 ����Ru�gk�eREV�!+��1�`���<S}�P�5C4O[T�ŅՔ`��

�ջ�'�Yp,-� ��F�Uy�di����0%���1�з�ex�^��F&���d{������aRcטėyy������h���se�1,�?+�E/�9�_E,f���~G��m&Y���ಧR���8���w�j
&yp���1 �W�?
�n�f%[Y�!�� �)Չ0����5]�N�z#x���.��{ox�c�b������}�5���m�W)��=/�3ۖ�?C�o����N�M���������db�U�WF-
���e$������e�K�
* L��s쎬C����/2�����C�P/�	�����X���A�8����}W�s�����"^{ldjT��[/&�C�&M�2�*A�i{��Mu}պ��x/]��U����_��KY��Ӵᴿ���%&]��,x���e�^�X���\L\��<���"��Lǥ���	�p�.�$F����P��~��]l`��bA��
.v}*,v�����9�oW�߂�*	A�(�����������&ǣ�@��i?jB% �S�]�i*���,���Xax�:8Y�	A�bY�����P�T ��?� � ��b�**4UF��РEp��M(�g�M�*0>�ųq	L�):�-q��L�V$���[<e�)#y�t��P��Ǯ�Z��?�Z�6ݞ�k�Dd�M6�g��d������
K�&CZY�����<oG/���áR!|�H�6q>c{�.�K*P��\�e��,��!�^'�u2�/g֢}�y���0##�t*�ى�H%1��0s�Vz���k@�qޕNr��ԸL(<~յ������Şt����;ȫ�u3Z&�e ���Ca?����0��!�����j�h��Hh�Y jv[��23�N=x�O�����Y�ZB�C�&�5��gP��{�����BNѽF~̄�Z§ 3sp��<�N?��G��d.m��:��AZ�fR�~����N � !����h�P#��K�C��wY4�.��v���r֧���X,�(�,�ϐqEb�݄���t��vʳO���	�{LD�iڪ�,ǋ�tS-�C&����:�ؓy����H{ߨW"` �:@��z2�8���k�;�����M�wI��*g�V�C5��E��	.����|��#Z�]��@����5�u����`/X�I ��q�"	y�������,�_�,U�{���j�j�_b4���CR��ޏ�F�SZ:I�rL�ܼ��H�>�9[8�]Ҵ�q�$��?�%O�S�b�Hj[���tJG�3P�uږnم`d�p̼�T���1�o0EB�~���G�\�&�n�|���GMT��6	�z������"�PMI��^^���B��J�s���跹#N8۹!ܸN ��s�*�==�N�`��Ì�b� �m�����׽/j�NZ#�x�8zy��1��V���<$�}૵�H�n��߽�q���y���t�F8��V��Yk�<q�Q|�!��#�&;p���Y\�MR�8!��.�"�|���i�s�ֶ�?��������л �E3`�ۙ�C������Θ���:Gq�v�^��t9�|�_�N����5��� �78�C�Ù}a������U3.厵��M Lʦ�<2��:�Ku4dM�'
�$,/��c$E���v����%j,�9�`9�<<`kp��&�:��$X|��}���P~<��F��8-X^ک@���eh���ӫ|�����,���7�|v��Xln�s�)�C�h�b�n�6ІT�Q͵O����.D ���h��A2��X�