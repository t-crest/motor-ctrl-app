-- DOC_Axis_Periphs_patmos.vhd

-- Generated using ACDS version 14.0 200 at 2015.08.07.09:58:31

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DOC_Axis_Periphs_patmos is
	port (
		drive0_adc_sync_dat_u           : in  std_logic                     := '0';             --              drive0_adc.sync_dat_u
		drive0_adc_sync_dat_w           : in  std_logic                     := '0';             --                        .sync_dat_w
		drive0_adc_overcurrent          : out std_logic;                                        --                        .overcurrent
		drive0_pwm_carrier              : out std_logic_vector(15 downto 0);                    --              drive0_pwm.carrier
		drive0_pwm_carrier_latch        : out std_logic;                                        --                        .carrier_latch
		drive0_pwm_encoder_strobe_n     : out std_logic;                                        --                        .encoder_strobe_n
		drive0_pwm_u_h                  : out std_logic;                                        --                        .u_h
		drive0_pwm_u_l                  : out std_logic;                                        --                        .u_l
		drive0_pwm_v_h                  : out std_logic;                                        --                        .v_h
		drive0_pwm_v_l                  : out std_logic;                                        --                        .v_l
		drive0_pwm_w_h                  : out std_logic;                                        --                        .w_h
		drive0_pwm_w_l                  : out std_logic;                                        --                        .w_l
		drive0_sm_overcurrent           : in  std_logic                     := '0';             --               drive0_sm.overcurrent
		drive0_sm_overvoltage           : in  std_logic                     := '0';             --                        .overvoltage
		drive0_sm_undervoltage          : in  std_logic                     := '0';             --                        .undervoltage
		drive0_sm_chopper               : in  std_logic                     := '0';             --                        .chopper
		drive0_sm_dc_link_clk_err       : in  std_logic                     := '0';             --                        .dc_link_clk_err
		drive0_sm_igbt_err              : in  std_logic                     := '0';             --                        .igbt_err
		drive0_sm_error_out             : out std_logic;                                        --                        .error_out
		drive0_sm_overcurrent_latch     : out std_logic;                                        --                        .overcurrent_latch
		drive0_sm_overvoltage_latch     : out std_logic;                                        --                        .overvoltage_latch
		drive0_sm_undervoltage_latch    : out std_logic;                                        --                        .undervoltage_latch
		drive0_sm_dc_link_clk_err_latch : out std_logic;                                        --                        .dc_link_clk_err_latch
		drive0_sm_igbt_err_latch        : out std_logic;                                        --                        .igbt_err_latch
		drive0_sm_chopper_latch         : out std_logic;                                        --                        .chopper_latch
		drive0_adc_pow_sync_dat_u       : in  std_logic                     := '0';             --          drive0_adc_pow.sync_dat_u
		drive0_adc_pow_sync_dat_w       : in  std_logic                     := '0';             --                        .sync_dat_w
		drive0_adc_pow_overcurrent      : out std_logic;                                        --                        .overcurrent
		clk_adc_in_clk                  : in  std_logic                     := '0';             --              clk_adc_in.clk
		drive0_biss_coe_ch1_MA          : out std_logic;                                        --             drive0_biss.coe_ch1_MA
		drive0_biss_coe_ch1_MO          : out std_logic;                                        --                        .coe_ch1_MO
		drive0_biss_coe_ch1_SL          : in  std_logic                     := '0';             --                        .coe_ch1_SL
		drive0_biss_coe_ch1_EOT         : out std_logic;                                        --                        .coe_ch1_EOT
		drive0_biss_get_sens            : in  std_logic                     := '0';             --                        .get_sens
		drive0_doc_pwm_sync_out_export  : out std_logic;                                        -- drive0_doc_pwm_sync_out.export
		drive0_doc_pwm_sync_in_export   : in  std_logic                     := '0';             --  drive0_doc_pwm_sync_in.export
		drive0_doc_adc_irq_irq          : out std_logic;                                        --      drive0_doc_adc_irq.irq
		drive0_doc_adc_pow_irq_irq      : out std_logic;                                        --  drive0_doc_adc_pow_irq.irq
		avs_periph_slave_waitrequest    : out std_logic;                                        --        avs_periph_slave.waitrequest
		avs_periph_slave_readdata       : out std_logic_vector(31 downto 0);                    --                        .readdata
		avs_periph_slave_readdatavalid  : out std_logic;                                        --                        .readdatavalid
		avs_periph_slave_burstcount     : in  std_logic_vector(0 downto 0)  := (others => '0'); --                        .burstcount
		avs_periph_slave_writedata      : in  std_logic_vector(31 downto 0) := (others => '0'); --                        .writedata
		avs_periph_slave_address        : in  std_logic_vector(11 downto 0) := (others => '0'); --                        .address
		avs_periph_slave_write          : in  std_logic                     := '0';             --                        .write
		avs_periph_slave_read           : in  std_logic                     := '0';             --                        .read
		avs_periph_slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => '0'); --                        .byteenable
		avs_periph_slave_debugaccess    : in  std_logic                     := '0';             --                        .debugaccess
		reset_reset_n                   : in  std_logic                     := '0';             --                   reset.reset_n
		clk_50_clk                      : in  std_logic                     := '0';             --                  clk_50.clk
		clk_80_clk                      : in  std_logic                     := '0';             --                  clk_80.clk
		reset_80_reset_n                : in  std_logic                     := '0'              --                reset_80.reset_n
	);
end entity DOC_Axis_Periphs_patmos;

architecture rtl of DOC_Axis_Periphs_patmos is
	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(11 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component DOC_Axis_Periphs_patmos_drive0 is
		port (
			clk_adc_clk               : in  std_logic                     := 'X';             -- clk
			reset_reset_n             : in  std_logic                     := 'X';             -- reset_n
			clk_periph_clk            : in  std_logic                     := 'X';             -- clk
			reset_periph_reset_n      : in  std_logic                     := 'X';             -- reset_n
			doc_adc_avs_write_n       : in  std_logic                     := 'X';             -- write_n
			doc_adc_avs_read_n        : in  std_logic                     := 'X';             -- read_n
			doc_adc_avs_address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			doc_adc_avs_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			doc_adc_avs_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			doc_adc_irq_irq           : out std_logic;                                        -- irq
			doc_pwm_avs_write_n       : in  std_logic                     := 'X';             -- write_n
			doc_pwm_avs_read_n        : in  std_logic                     := 'X';             -- read_n
			doc_pwm_avs_address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			doc_pwm_avs_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			doc_pwm_avs_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			doc_sm_avs_write_n        : in  std_logic                     := 'X';             -- write_n
			doc_sm_avs_read_n         : in  std_logic                     := 'X';             -- read_n
			doc_sm_avs_address        : in  std_logic                     := 'X';             -- address
			doc_sm_avs_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			doc_sm_avs_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			doc_adc_pow_avs_write_n   : in  std_logic                     := 'X';             -- write_n
			doc_adc_pow_avs_read_n    : in  std_logic                     := 'X';             -- read_n
			doc_adc_pow_avs_address   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			doc_adc_pow_avs_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			doc_adc_pow_avs_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			doc_adc_pow_irq_irq       : out std_logic;                                        -- irq
			doc_pwm_sync_out_export   : out std_logic;                                        -- export
			doc_pwm_sync_in_export    : in  std_logic                     := 'X';             -- export
			adc_pow_sync_dat_u        : in  std_logic                     := 'X';             -- sync_dat_u
			adc_pow_sync_dat_w        : in  std_logic                     := 'X';             -- sync_dat_w
			adc_pow_overcurrent       : out std_logic;                                        -- overcurrent
			adc_sync_dat_u            : in  std_logic                     := 'X';             -- sync_dat_u
			adc_sync_dat_w            : in  std_logic                     := 'X';             -- sync_dat_w
			adc_overcurrent           : out std_logic;                                        -- overcurrent
			pwm_carrier               : out std_logic_vector(15 downto 0);                    -- carrier
			pwm_carrier_latch         : out std_logic;                                        -- carrier_latch
			pwm_encoder_strobe_n      : out std_logic;                                        -- encoder_strobe_n
			pwm_u_h                   : out std_logic;                                        -- u_h
			pwm_u_l                   : out std_logic;                                        -- u_l
			pwm_v_h                   : out std_logic;                                        -- v_h
			pwm_v_l                   : out std_logic;                                        -- v_l
			pwm_w_h                   : out std_logic;                                        -- w_h
			pwm_w_l                   : out std_logic;                                        -- w_l
			sm_overcurrent            : in  std_logic                     := 'X';             -- overcurrent
			sm_overvoltage            : in  std_logic                     := 'X';             -- overvoltage
			sm_undervoltage           : in  std_logic                     := 'X';             -- undervoltage
			sm_chopper                : in  std_logic                     := 'X';             -- chopper
			sm_dc_link_clk_err        : in  std_logic                     := 'X';             -- dc_link_clk_err
			sm_igbt_err               : in  std_logic                     := 'X';             -- igbt_err
			sm_error_out              : out std_logic;                                        -- error_out
			sm_overcurrent_latch      : out std_logic;                                        -- overcurrent_latch
			sm_overvoltage_latch      : out std_logic;                                        -- overvoltage_latch
			sm_undervoltage_latch     : out std_logic;                                        -- undervoltage_latch
			sm_dc_link_clk_err_latch  : out std_logic;                                        -- dc_link_clk_err_latch
			sm_igbt_err_latch         : out std_logic;                                        -- igbt_err_latch
			sm_chopper_latch          : out std_logic;                                        -- chopper_latch
			doc_biss_avs_write_n      : in  std_logic                     := 'X';             -- write_n
			doc_biss_avs_read_n       : in  std_logic                     := 'X';             -- read_n
			doc_biss_avs_address      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			doc_biss_avs_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			doc_biss_avs_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			doc_biss_avs_chipselect_n : in  std_logic                     := 'X';             -- chipselect_n
			doc_biss_coe_ch1_MA       : out std_logic;                                        -- coe_ch1_MA
			doc_biss_coe_ch1_MO       : out std_logic;                                        -- coe_ch1_MO
			doc_biss_coe_ch1_SL       : in  std_logic                     := 'X';             -- coe_ch1_SL
			doc_biss_coe_ch1_EOT      : out std_logic;                                        -- coe_ch1_EOT
			doc_biss_get_sens         : in  std_logic                     := 'X';             -- get_sens
			doc_biss_irq_irq          : out std_logic                                         -- irq
		);
	end component DOC_Axis_Periphs_patmos_drive0;

	component DOC_Axis_Periphs_patmos_mm_interconnect_0 is
		port (
			clk_int_50_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			clock_crossing_m0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			drive0_reset_periph_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			clock_crossing_m0_address                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clock_crossing_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			clock_crossing_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			clock_crossing_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock_crossing_m0_read                              : in  std_logic                     := 'X';             -- read
			clock_crossing_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			clock_crossing_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			clock_crossing_m0_write                             : in  std_logic                     := 'X';             -- write
			clock_crossing_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_crossing_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			drive0_doc_adc_avs_address                          : out std_logic_vector(3 downto 0);                     -- address
			drive0_doc_adc_avs_write                            : out std_logic;                                        -- write
			drive0_doc_adc_avs_read                             : out std_logic;                                        -- read
			drive0_doc_adc_avs_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			drive0_doc_adc_avs_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			drive0_doc_adc_pow_avs_address                      : out std_logic_vector(3 downto 0);                     -- address
			drive0_doc_adc_pow_avs_write                        : out std_logic;                                        -- write
			drive0_doc_adc_pow_avs_read                         : out std_logic;                                        -- read
			drive0_doc_adc_pow_avs_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			drive0_doc_adc_pow_avs_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			drive0_doc_biss_avs_address                         : out std_logic_vector(5 downto 0);                     -- address
			drive0_doc_biss_avs_write                           : out std_logic;                                        -- write
			drive0_doc_biss_avs_read                            : out std_logic;                                        -- read
			drive0_doc_biss_avs_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			drive0_doc_biss_avs_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			drive0_doc_biss_avs_chipselect                      : out std_logic;                                        -- chipselect
			drive0_doc_pwm_avs_address                          : out std_logic_vector(3 downto 0);                     -- address
			drive0_doc_pwm_avs_write                            : out std_logic;                                        -- write
			drive0_doc_pwm_avs_read                             : out std_logic;                                        -- read
			drive0_doc_pwm_avs_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			drive0_doc_pwm_avs_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			drive0_doc_sm_avs_address                           : out std_logic_vector(0 downto 0);                     -- address
			drive0_doc_sm_avs_write                             : out std_logic;                                        -- write
			drive0_doc_sm_avs_read                              : out std_logic;                                        -- read
			drive0_doc_sm_avs_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			drive0_doc_sm_avs_writedata                         : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component DOC_Axis_Periphs_patmos_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal clock_crossing_m0_burstcount                               : std_logic_vector(0 downto 0);  -- clock_crossing:m0_burstcount -> mm_interconnect_0:clock_crossing_m0_burstcount
	signal clock_crossing_m0_waitrequest                              : std_logic;                     -- mm_interconnect_0:clock_crossing_m0_waitrequest -> clock_crossing:m0_waitrequest
	signal clock_crossing_m0_address                                  : std_logic_vector(11 downto 0); -- clock_crossing:m0_address -> mm_interconnect_0:clock_crossing_m0_address
	signal clock_crossing_m0_writedata                                : std_logic_vector(31 downto 0); -- clock_crossing:m0_writedata -> mm_interconnect_0:clock_crossing_m0_writedata
	signal clock_crossing_m0_write                                    : std_logic;                     -- clock_crossing:m0_write -> mm_interconnect_0:clock_crossing_m0_write
	signal clock_crossing_m0_read                                     : std_logic;                     -- clock_crossing:m0_read -> mm_interconnect_0:clock_crossing_m0_read
	signal clock_crossing_m0_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:clock_crossing_m0_readdata -> clock_crossing:m0_readdata
	signal clock_crossing_m0_debugaccess                              : std_logic;                     -- clock_crossing:m0_debugaccess -> mm_interconnect_0:clock_crossing_m0_debugaccess
	signal clock_crossing_m0_byteenable                               : std_logic_vector(3 downto 0);  -- clock_crossing:m0_byteenable -> mm_interconnect_0:clock_crossing_m0_byteenable
	signal clock_crossing_m0_readdatavalid                            : std_logic;                     -- mm_interconnect_0:clock_crossing_m0_readdatavalid -> clock_crossing:m0_readdatavalid
	signal mm_interconnect_0_drive0_doc_pwm_avs_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:drive0_doc_pwm_avs_writedata -> drive0:doc_pwm_avs_writedata
	signal mm_interconnect_0_drive0_doc_pwm_avs_address               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:drive0_doc_pwm_avs_address -> drive0:doc_pwm_avs_address
	signal mm_interconnect_0_drive0_doc_pwm_avs_write                 : std_logic;                     -- mm_interconnect_0:drive0_doc_pwm_avs_write -> mm_interconnect_0_drive0_doc_pwm_avs_write:in
	signal mm_interconnect_0_drive0_doc_pwm_avs_read                  : std_logic;                     -- mm_interconnect_0:drive0_doc_pwm_avs_read -> mm_interconnect_0_drive0_doc_pwm_avs_read:in
	signal mm_interconnect_0_drive0_doc_pwm_avs_readdata              : std_logic_vector(31 downto 0); -- drive0:doc_pwm_avs_readdata -> mm_interconnect_0:drive0_doc_pwm_avs_readdata
	signal mm_interconnect_0_drive0_doc_sm_avs_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:drive0_doc_sm_avs_writedata -> drive0:doc_sm_avs_writedata
	signal mm_interconnect_0_drive0_doc_sm_avs_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:drive0_doc_sm_avs_address -> drive0:doc_sm_avs_address
	signal mm_interconnect_0_drive0_doc_sm_avs_write                  : std_logic;                     -- mm_interconnect_0:drive0_doc_sm_avs_write -> mm_interconnect_0_drive0_doc_sm_avs_write:in
	signal mm_interconnect_0_drive0_doc_sm_avs_read                   : std_logic;                     -- mm_interconnect_0:drive0_doc_sm_avs_read -> mm_interconnect_0_drive0_doc_sm_avs_read:in
	signal mm_interconnect_0_drive0_doc_sm_avs_readdata               : std_logic_vector(31 downto 0); -- drive0:doc_sm_avs_readdata -> mm_interconnect_0:drive0_doc_sm_avs_readdata
	signal mm_interconnect_0_drive0_doc_adc_avs_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:drive0_doc_adc_avs_writedata -> drive0:doc_adc_avs_writedata
	signal mm_interconnect_0_drive0_doc_adc_avs_address               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:drive0_doc_adc_avs_address -> drive0:doc_adc_avs_address
	signal mm_interconnect_0_drive0_doc_adc_avs_write                 : std_logic;                     -- mm_interconnect_0:drive0_doc_adc_avs_write -> mm_interconnect_0_drive0_doc_adc_avs_write:in
	signal mm_interconnect_0_drive0_doc_adc_avs_read                  : std_logic;                     -- mm_interconnect_0:drive0_doc_adc_avs_read -> mm_interconnect_0_drive0_doc_adc_avs_read:in
	signal mm_interconnect_0_drive0_doc_adc_avs_readdata              : std_logic_vector(31 downto 0); -- drive0:doc_adc_avs_readdata -> mm_interconnect_0:drive0_doc_adc_avs_readdata
	signal mm_interconnect_0_drive0_doc_adc_pow_avs_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:drive0_doc_adc_pow_avs_writedata -> drive0:doc_adc_pow_avs_writedata
	signal mm_interconnect_0_drive0_doc_adc_pow_avs_address           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:drive0_doc_adc_pow_avs_address -> drive0:doc_adc_pow_avs_address
	signal mm_interconnect_0_drive0_doc_adc_pow_avs_write             : std_logic;                     -- mm_interconnect_0:drive0_doc_adc_pow_avs_write -> mm_interconnect_0_drive0_doc_adc_pow_avs_write:in
	signal mm_interconnect_0_drive0_doc_adc_pow_avs_read              : std_logic;                     -- mm_interconnect_0:drive0_doc_adc_pow_avs_read -> mm_interconnect_0_drive0_doc_adc_pow_avs_read:in
	signal mm_interconnect_0_drive0_doc_adc_pow_avs_readdata          : std_logic_vector(31 downto 0); -- drive0:doc_adc_pow_avs_readdata -> mm_interconnect_0:drive0_doc_adc_pow_avs_readdata
	signal mm_interconnect_0_drive0_doc_biss_avs_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:drive0_doc_biss_avs_writedata -> drive0:doc_biss_avs_writedata
	signal mm_interconnect_0_drive0_doc_biss_avs_address              : std_logic_vector(5 downto 0);  -- mm_interconnect_0:drive0_doc_biss_avs_address -> drive0:doc_biss_avs_address
	signal mm_interconnect_0_drive0_doc_biss_avs_chipselect           : std_logic;                     -- mm_interconnect_0:drive0_doc_biss_avs_chipselect -> mm_interconnect_0_drive0_doc_biss_avs_chipselect:in
	signal mm_interconnect_0_drive0_doc_biss_avs_write                : std_logic;                     -- mm_interconnect_0:drive0_doc_biss_avs_write -> mm_interconnect_0_drive0_doc_biss_avs_write:in
	signal mm_interconnect_0_drive0_doc_biss_avs_read                 : std_logic;                     -- mm_interconnect_0:drive0_doc_biss_avs_read -> mm_interconnect_0_drive0_doc_biss_avs_read:in
	signal mm_interconnect_0_drive0_doc_biss_avs_readdata             : std_logic_vector(31 downto 0); -- drive0:doc_biss_avs_readdata -> mm_interconnect_0:drive0_doc_biss_avs_readdata
	signal rst_controller_reset_out_reset                             : std_logic;                     -- rst_controller:reset_out -> [clock_crossing:m0_reset, mm_interconnect_0:clock_crossing_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:drive0_reset_periph_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                         : std_logic;                     -- rst_controller_001:reset_out -> clock_crossing:s0_reset
	signal reset_reset_n_ports_inv                                    : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal reset_80_reset_n_ports_inv                                 : std_logic;                     -- reset_80_reset_n:inv -> rst_controller_001:reset_in0
	signal mm_interconnect_0_drive0_doc_pwm_avs_write_ports_inv       : std_logic;                     -- mm_interconnect_0_drive0_doc_pwm_avs_write:inv -> drive0:doc_pwm_avs_write_n
	signal mm_interconnect_0_drive0_doc_pwm_avs_read_ports_inv        : std_logic;                     -- mm_interconnect_0_drive0_doc_pwm_avs_read:inv -> drive0:doc_pwm_avs_read_n
	signal mm_interconnect_0_drive0_doc_sm_avs_write_ports_inv        : std_logic;                     -- mm_interconnect_0_drive0_doc_sm_avs_write:inv -> drive0:doc_sm_avs_write_n
	signal mm_interconnect_0_drive0_doc_sm_avs_read_ports_inv         : std_logic;                     -- mm_interconnect_0_drive0_doc_sm_avs_read:inv -> drive0:doc_sm_avs_read_n
	signal mm_interconnect_0_drive0_doc_adc_avs_write_ports_inv       : std_logic;                     -- mm_interconnect_0_drive0_doc_adc_avs_write:inv -> drive0:doc_adc_avs_write_n
	signal mm_interconnect_0_drive0_doc_adc_avs_read_ports_inv        : std_logic;                     -- mm_interconnect_0_drive0_doc_adc_avs_read:inv -> drive0:doc_adc_avs_read_n
	signal mm_interconnect_0_drive0_doc_adc_pow_avs_write_ports_inv   : std_logic;                     -- mm_interconnect_0_drive0_doc_adc_pow_avs_write:inv -> drive0:doc_adc_pow_avs_write_n
	signal mm_interconnect_0_drive0_doc_adc_pow_avs_read_ports_inv    : std_logic;                     -- mm_interconnect_0_drive0_doc_adc_pow_avs_read:inv -> drive0:doc_adc_pow_avs_read_n
	signal mm_interconnect_0_drive0_doc_biss_avs_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_drive0_doc_biss_avs_chipselect:inv -> drive0:doc_biss_avs_chipselect_n
	signal mm_interconnect_0_drive0_doc_biss_avs_write_ports_inv      : std_logic;                     -- mm_interconnect_0_drive0_doc_biss_avs_write:inv -> drive0:doc_biss_avs_write_n
	signal mm_interconnect_0_drive0_doc_biss_avs_read_ports_inv       : std_logic;                     -- mm_interconnect_0_drive0_doc_biss_avs_read:inv -> drive0:doc_biss_avs_read_n

begin

	clock_crossing : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 12,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 2,
			RESPONSE_FIFO_DEPTH => 2,
			MASTER_SYNC_DEPTH   => 3,
			SLAVE_SYNC_DEPTH    => 3
		)
		port map (
			m0_clk           => clk_50_clk,                         --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,     -- m0_reset.reset
			s0_clk           => clk_80_clk,                         --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset, -- s0_reset.reset
			s0_waitrequest   => avs_periph_slave_waitrequest,       --       s0.waitrequest
			s0_readdata      => avs_periph_slave_readdata,          --         .readdata
			s0_readdatavalid => avs_periph_slave_readdatavalid,     --         .readdatavalid
			s0_burstcount    => avs_periph_slave_burstcount,        --         .burstcount
			s0_writedata     => avs_periph_slave_writedata,         --         .writedata
			s0_address       => avs_periph_slave_address,           --         .address
			s0_write         => avs_periph_slave_write,             --         .write
			s0_read          => avs_periph_slave_read,              --         .read
			s0_byteenable    => avs_periph_slave_byteenable,        --         .byteenable
			s0_debugaccess   => avs_periph_slave_debugaccess,       --         .debugaccess
			m0_waitrequest   => clock_crossing_m0_waitrequest,      --       m0.waitrequest
			m0_readdata      => clock_crossing_m0_readdata,         --         .readdata
			m0_readdatavalid => clock_crossing_m0_readdatavalid,    --         .readdatavalid
			m0_burstcount    => clock_crossing_m0_burstcount,       --         .burstcount
			m0_writedata     => clock_crossing_m0_writedata,        --         .writedata
			m0_address       => clock_crossing_m0_address,          --         .address
			m0_write         => clock_crossing_m0_write,            --         .write
			m0_read          => clock_crossing_m0_read,             --         .read
			m0_byteenable    => clock_crossing_m0_byteenable,       --         .byteenable
			m0_debugaccess   => clock_crossing_m0_debugaccess       --         .debugaccess
		);

	drive0 : component DOC_Axis_Periphs_patmos_drive0
		port map (
			clk_adc_clk               => clk_adc_in_clk,                                             --          clk_adc.clk
			reset_reset_n             => reset_reset_n,                                              --            reset.reset_n
			clk_periph_clk            => clk_50_clk,                                                 --       clk_periph.clk
			reset_periph_reset_n      => reset_reset_n,                                              --     reset_periph.reset_n
			doc_adc_avs_write_n       => mm_interconnect_0_drive0_doc_adc_avs_write_ports_inv,       --      doc_adc_avs.write_n
			doc_adc_avs_read_n        => mm_interconnect_0_drive0_doc_adc_avs_read_ports_inv,        --                 .read_n
			doc_adc_avs_address       => mm_interconnect_0_drive0_doc_adc_avs_address,               --                 .address
			doc_adc_avs_writedata     => mm_interconnect_0_drive0_doc_adc_avs_writedata,             --                 .writedata
			doc_adc_avs_readdata      => mm_interconnect_0_drive0_doc_adc_avs_readdata,              --                 .readdata
			doc_adc_irq_irq           => drive0_doc_adc_irq_irq,                                     --      doc_adc_irq.irq
			doc_pwm_avs_write_n       => mm_interconnect_0_drive0_doc_pwm_avs_write_ports_inv,       --      doc_pwm_avs.write_n
			doc_pwm_avs_read_n        => mm_interconnect_0_drive0_doc_pwm_avs_read_ports_inv,        --                 .read_n
			doc_pwm_avs_address       => mm_interconnect_0_drive0_doc_pwm_avs_address,               --                 .address
			doc_pwm_avs_writedata     => mm_interconnect_0_drive0_doc_pwm_avs_writedata,             --                 .writedata
			doc_pwm_avs_readdata      => mm_interconnect_0_drive0_doc_pwm_avs_readdata,              --                 .readdata
			doc_sm_avs_write_n        => mm_interconnect_0_drive0_doc_sm_avs_write_ports_inv,        --       doc_sm_avs.write_n
			doc_sm_avs_read_n         => mm_interconnect_0_drive0_doc_sm_avs_read_ports_inv,         --                 .read_n
			doc_sm_avs_address        => mm_interconnect_0_drive0_doc_sm_avs_address(0),             --                 .address
			doc_sm_avs_writedata      => mm_interconnect_0_drive0_doc_sm_avs_writedata,              --                 .writedata
			doc_sm_avs_readdata       => mm_interconnect_0_drive0_doc_sm_avs_readdata,               --                 .readdata
			doc_adc_pow_avs_write_n   => mm_interconnect_0_drive0_doc_adc_pow_avs_write_ports_inv,   --  doc_adc_pow_avs.write_n
			doc_adc_pow_avs_read_n    => mm_interconnect_0_drive0_doc_adc_pow_avs_read_ports_inv,    --                 .read_n
			doc_adc_pow_avs_address   => mm_interconnect_0_drive0_doc_adc_pow_avs_address,           --                 .address
			doc_adc_pow_avs_writedata => mm_interconnect_0_drive0_doc_adc_pow_avs_writedata,         --                 .writedata
			doc_adc_pow_avs_readdata  => mm_interconnect_0_drive0_doc_adc_pow_avs_readdata,          --                 .readdata
			doc_adc_pow_irq_irq       => drive0_doc_adc_pow_irq_irq,                                 --  doc_adc_pow_irq.irq
			doc_pwm_sync_out_export   => drive0_doc_pwm_sync_out_export,                             -- doc_pwm_sync_out.export
			doc_pwm_sync_in_export    => drive0_doc_pwm_sync_in_export,                              --  doc_pwm_sync_in.export
			adc_pow_sync_dat_u        => drive0_adc_pow_sync_dat_u,                                  --          adc_pow.sync_dat_u
			adc_pow_sync_dat_w        => drive0_adc_pow_sync_dat_w,                                  --                 .sync_dat_w
			adc_pow_overcurrent       => drive0_adc_pow_overcurrent,                                 --                 .overcurrent
			adc_sync_dat_u            => drive0_adc_sync_dat_u,                                      --              adc.sync_dat_u
			adc_sync_dat_w            => drive0_adc_sync_dat_w,                                      --                 .sync_dat_w
			adc_overcurrent           => drive0_adc_overcurrent,                                     --                 .overcurrent
			pwm_carrier               => drive0_pwm_carrier,                                         --              pwm.carrier
			pwm_carrier_latch         => drive0_pwm_carrier_latch,                                   --                 .carrier_latch
			pwm_encoder_strobe_n      => drive0_pwm_encoder_strobe_n,                                --                 .encoder_strobe_n
			pwm_u_h                   => drive0_pwm_u_h,                                             --                 .u_h
			pwm_u_l                   => drive0_pwm_u_l,                                             --                 .u_l
			pwm_v_h                   => drive0_pwm_v_h,                                             --                 .v_h
			pwm_v_l                   => drive0_pwm_v_l,                                             --                 .v_l
			pwm_w_h                   => drive0_pwm_w_h,                                             --                 .w_h
			pwm_w_l                   => drive0_pwm_w_l,                                             --                 .w_l
			sm_overcurrent            => drive0_sm_overcurrent,                                      --               sm.overcurrent
			sm_overvoltage            => drive0_sm_overvoltage,                                      --                 .overvoltage
			sm_undervoltage           => drive0_sm_undervoltage,                                     --                 .undervoltage
			sm_chopper                => drive0_sm_chopper,                                          --                 .chopper
			sm_dc_link_clk_err        => drive0_sm_dc_link_clk_err,                                  --                 .dc_link_clk_err
			sm_igbt_err               => drive0_sm_igbt_err,                                         --                 .igbt_err
			sm_error_out              => drive0_sm_error_out,                                        --                 .error_out
			sm_overcurrent_latch      => drive0_sm_overcurrent_latch,                                --                 .overcurrent_latch
			sm_overvoltage_latch      => drive0_sm_overvoltage_latch,                                --                 .overvoltage_latch
			sm_undervoltage_latch     => drive0_sm_undervoltage_latch,                               --                 .undervoltage_latch
			sm_dc_link_clk_err_latch  => drive0_sm_dc_link_clk_err_latch,                            --                 .dc_link_clk_err_latch
			sm_igbt_err_latch         => drive0_sm_igbt_err_latch,                                   --                 .igbt_err_latch
			sm_chopper_latch          => drive0_sm_chopper_latch,                                    --                 .chopper_latch
			doc_biss_avs_write_n      => mm_interconnect_0_drive0_doc_biss_avs_write_ports_inv,      --     doc_biss_avs.write_n
			doc_biss_avs_read_n       => mm_interconnect_0_drive0_doc_biss_avs_read_ports_inv,       --                 .read_n
			doc_biss_avs_address      => mm_interconnect_0_drive0_doc_biss_avs_address,              --                 .address
			doc_biss_avs_writedata    => mm_interconnect_0_drive0_doc_biss_avs_writedata,            --                 .writedata
			doc_biss_avs_readdata     => mm_interconnect_0_drive0_doc_biss_avs_readdata,             --                 .readdata
			doc_biss_avs_chipselect_n => mm_interconnect_0_drive0_doc_biss_avs_chipselect_ports_inv, --                 .chipselect_n
			doc_biss_coe_ch1_MA       => drive0_biss_coe_ch1_MA,                                     --         doc_biss.coe_ch1_MA
			doc_biss_coe_ch1_MO       => drive0_biss_coe_ch1_MO,                                     --                 .coe_ch1_MO
			doc_biss_coe_ch1_SL       => drive0_biss_coe_ch1_SL,                                     --                 .coe_ch1_SL
			doc_biss_coe_ch1_EOT      => drive0_biss_coe_ch1_EOT,                                    --                 .coe_ch1_EOT
			doc_biss_get_sens         => drive0_biss_get_sens,                                       --                 .get_sens
			doc_biss_irq_irq          => open                                                        --     doc_biss_irq.irq
		);

	mm_interconnect_0 : component DOC_Axis_Periphs_patmos_mm_interconnect_0
		port map (
			clk_int_50_clk_clk                                  => clk_50_clk,                                         --                                clk_int_50_clk.clk
			clock_crossing_m0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                     -- clock_crossing_m0_reset_reset_bridge_in_reset.reset
			drive0_reset_periph_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                     --     drive0_reset_periph_reset_bridge_in_reset.reset
			clock_crossing_m0_address                           => clock_crossing_m0_address,                          --                             clock_crossing_m0.address
			clock_crossing_m0_waitrequest                       => clock_crossing_m0_waitrequest,                      --                                              .waitrequest
			clock_crossing_m0_burstcount                        => clock_crossing_m0_burstcount,                       --                                              .burstcount
			clock_crossing_m0_byteenable                        => clock_crossing_m0_byteenable,                       --                                              .byteenable
			clock_crossing_m0_read                              => clock_crossing_m0_read,                             --                                              .read
			clock_crossing_m0_readdata                          => clock_crossing_m0_readdata,                         --                                              .readdata
			clock_crossing_m0_readdatavalid                     => clock_crossing_m0_readdatavalid,                    --                                              .readdatavalid
			clock_crossing_m0_write                             => clock_crossing_m0_write,                            --                                              .write
			clock_crossing_m0_writedata                         => clock_crossing_m0_writedata,                        --                                              .writedata
			clock_crossing_m0_debugaccess                       => clock_crossing_m0_debugaccess,                      --                                              .debugaccess
			drive0_doc_adc_avs_address                          => mm_interconnect_0_drive0_doc_adc_avs_address,       --                            drive0_doc_adc_avs.address
			drive0_doc_adc_avs_write                            => mm_interconnect_0_drive0_doc_adc_avs_write,         --                                              .write
			drive0_doc_adc_avs_read                             => mm_interconnect_0_drive0_doc_adc_avs_read,          --                                              .read
			drive0_doc_adc_avs_readdata                         => mm_interconnect_0_drive0_doc_adc_avs_readdata,      --                                              .readdata
			drive0_doc_adc_avs_writedata                        => mm_interconnect_0_drive0_doc_adc_avs_writedata,     --                                              .writedata
			drive0_doc_adc_pow_avs_address                      => mm_interconnect_0_drive0_doc_adc_pow_avs_address,   --                        drive0_doc_adc_pow_avs.address
			drive0_doc_adc_pow_avs_write                        => mm_interconnect_0_drive0_doc_adc_pow_avs_write,     --                                              .write
			drive0_doc_adc_pow_avs_read                         => mm_interconnect_0_drive0_doc_adc_pow_avs_read,      --                                              .read
			drive0_doc_adc_pow_avs_readdata                     => mm_interconnect_0_drive0_doc_adc_pow_avs_readdata,  --                                              .readdata
			drive0_doc_adc_pow_avs_writedata                    => mm_interconnect_0_drive0_doc_adc_pow_avs_writedata, --                                              .writedata
			drive0_doc_biss_avs_address                         => mm_interconnect_0_drive0_doc_biss_avs_address,      --                           drive0_doc_biss_avs.address
			drive0_doc_biss_avs_write                           => mm_interconnect_0_drive0_doc_biss_avs_write,        --                                              .write
			drive0_doc_biss_avs_read                            => mm_interconnect_0_drive0_doc_biss_avs_read,         --                                              .read
			drive0_doc_biss_avs_readdata                        => mm_interconnect_0_drive0_doc_biss_avs_readdata,     --                                              .readdata
			drive0_doc_biss_avs_writedata                       => mm_interconnect_0_drive0_doc_biss_avs_writedata,    --                                              .writedata
			drive0_doc_biss_avs_chipselect                      => mm_interconnect_0_drive0_doc_biss_avs_chipselect,   --                                              .chipselect
			drive0_doc_pwm_avs_address                          => mm_interconnect_0_drive0_doc_pwm_avs_address,       --                            drive0_doc_pwm_avs.address
			drive0_doc_pwm_avs_write                            => mm_interconnect_0_drive0_doc_pwm_avs_write,         --                                              .write
			drive0_doc_pwm_avs_read                             => mm_interconnect_0_drive0_doc_pwm_avs_read,          --                                              .read
			drive0_doc_pwm_avs_readdata                         => mm_interconnect_0_drive0_doc_pwm_avs_readdata,      --                                              .readdata
			drive0_doc_pwm_avs_writedata                        => mm_interconnect_0_drive0_doc_pwm_avs_writedata,     --                                              .writedata
			drive0_doc_sm_avs_address                           => mm_interconnect_0_drive0_doc_sm_avs_address,        --                             drive0_doc_sm_avs.address
			drive0_doc_sm_avs_write                             => mm_interconnect_0_drive0_doc_sm_avs_write,          --                                              .write
			drive0_doc_sm_avs_read                              => mm_interconnect_0_drive0_doc_sm_avs_read,           --                                              .read
			drive0_doc_sm_avs_readdata                          => mm_interconnect_0_drive0_doc_sm_avs_readdata,       --                                              .readdata
			drive0_doc_sm_avs_writedata                         => mm_interconnect_0_drive0_doc_sm_avs_writedata       --                                              .writedata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_50_clk,                     --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_80_reset_n_ports_inv,         -- reset_in0.reset
			clk            => clk_80_clk,                         --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	reset_80_reset_n_ports_inv <= not reset_80_reset_n;

	mm_interconnect_0_drive0_doc_pwm_avs_write_ports_inv <= not mm_interconnect_0_drive0_doc_pwm_avs_write;

	mm_interconnect_0_drive0_doc_pwm_avs_read_ports_inv <= not mm_interconnect_0_drive0_doc_pwm_avs_read;

	mm_interconnect_0_drive0_doc_sm_avs_write_ports_inv <= not mm_interconnect_0_drive0_doc_sm_avs_write;

	mm_interconnect_0_drive0_doc_sm_avs_read_ports_inv <= not mm_interconnect_0_drive0_doc_sm_avs_read;

	mm_interconnect_0_drive0_doc_adc_avs_write_ports_inv <= not mm_interconnect_0_drive0_doc_adc_avs_write;

	mm_interconnect_0_drive0_doc_adc_avs_read_ports_inv <= not mm_interconnect_0_drive0_doc_adc_avs_read;

	mm_interconnect_0_drive0_doc_adc_pow_avs_write_ports_inv <= not mm_interconnect_0_drive0_doc_adc_pow_avs_write;

	mm_interconnect_0_drive0_doc_adc_pow_avs_read_ports_inv <= not mm_interconnect_0_drive0_doc_adc_pow_avs_read;

	mm_interconnect_0_drive0_doc_biss_avs_chipselect_ports_inv <= not mm_interconnect_0_drive0_doc_biss_avs_chipselect;

	mm_interconnect_0_drive0_doc_biss_avs_write_ports_inv <= not mm_interconnect_0_drive0_doc_biss_avs_write;

	mm_interconnect_0_drive0_doc_biss_avs_read_ports_inv <= not mm_interconnect_0_drive0_doc_biss_avs_read;

end architecture rtl; -- of DOC_Axis_Periphs_patmos
