��/  h$�p�̦[�)t��ׅ����^N_��?H4�ӝe2L�B���)k%���C&�)Fy���*�9�srq�},��(��z�I�e�A���_�.$�P����P�T�i4��:]+u�;�i�B|��yOܲF�L�ߖ�>�Y��#��L��"aQ��0�͵�9���K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<�P�����P��v͹	�$��)zuVB뼵=�~h]o
����-����%,@�`ٳ��K����\�zg�tݼ��%x.妀T��4] ���4^2$3I<N��褗���FR��L��B>SY�;��}���Zı�<%��3�OT�@EnPݣSW��*�C}XY������9?ƍ�t��L����!�"�.�[�,�WK���.�A�w��.o����6E�lW;M�)j>���/�����������>�)���A91���a��jk\��x?#q�iw0�@�r�X	�_D�j�������>+>��;}�ZJ��Q�RB�#c�z�i���$�e~cV�F�oF� �eS�����%�b�5�L�{c} �L��CAN�XC��g��X��_��G�z��]v��wp��<[�������u�fIC1�D��P9���%+��,��qЅ���M"��5K�F� �_�vj�`�Y��8넔y�(�=�\W���	�tZC�Y<�/�Bt�b��o8�6�Z�t�]�SV�VA4�g�OH�"
O��{����ٸ|񗿤,tIr�s��+���V�B[�4~:4[�h"��6Ul,ǀ��,s�`�D����,�s36	,�X�R���Ej�w�T��]��x����!�6q��Y[E
��3�Oi/#�"�z�\A����O�J�Te���2�~m���h�MN�~f��s4W�����ݭ3*��6�?R,Y�#�l$E�Uy������*F������.��v�K����a=,��7&��a]��s\a\�Iͩ#�o���*�����r��~�Pk��:��K
e��^����n`�a���}��W�L�P�]��~¡����=*+K��c�����d!�^HY��Ҿ�RKZ�6ıs��w
}E.�?��0@W�����D[�`���[�5�-�y|R����=��{F����$�����¯~geZx��2������o�o+J����D.�ݦO�@P���a��,5Q�9��b�͟���hg9i�������!��
$����Q��,?���x9Y�3 �m�4�BP(�yN^1ѽ�P����aM����k8y�z$;��Q��ߞ��f/\�/6��;��Z�p6N��7Q�6��4.�[~�P�*�&Q�]��\Y��d�q9v�5�*:b*I��s=����S����rӡN�"48ց��5������ZT��x��sJgAUg�d��]U�=���E���=���G����ej,g9��\ý�$��yx9�dm�����S*��M����Ϙ���B-�g�˃ �"^���K�1�4"i$R�$`������g�s]�&Zʓ� ��]8³&�Y*HH�fB����jTNI 2u6��-�l!R�"�� �*��uǖ��p�[��H�?����z�0�ř��տ3y*i������x'U��W�PE�0��;���B �n-�F��_X+�L�~w�j�����L����K�S�1���d� Y��%����{��K��)��,�F�3x���y���P��-���2�6��_���mب���,��j��G��iD�f�e��~??��©���XT���2P��J��=
��s� o�L*����Oj��� gӦ��]l��_��!<}�E�B�bo��X�W�[�Le=��a��8a�:�V���5��6+{\.!��%�+���DJ���wx�$������PR���`CW��xM�o�{\O����*~�O"���3wi�i��th�����^�d&����i����GB�S�,z:�[i*��ĕ��*>IqH��&z�A�oB��%gΒ�ƅ$�%il��$�~A���O� �R�0��ҹ�IR�x�ZiZa֚���n�ꈋ���V��f���cK~�4�l��u_� �@'��n?�#p�)b�v��	0nEd��y���!�L:� #�j+'Ӌ��/�۪��i�� R�) +��$�o�����ؿA�qȂ�����b���*N�AM:ʄc ��0��p��O�q���6��J<�.-�A�Q�Z�16<��rK_I�rm�F!���$��f��##/F��ߘ��8��.��D@���B�d��X�3�`k:�$[F6��ƯUO���=I��UL iYP��������'���p���_�h�K��QA!h��=T����w�gQ`]j3P�H�d�E�{R��.+�u��:7V��;^�A��8�0�qW#�Uo��6�4���ߞk�;�$�ƶ�#�*�Y�n?�̘�����f�(T�ߗ'���A_��S�B'���h��25����I�8�y'J1���Ә�h)�~wu:E�J!-���y�Vh�Q͟�Z�Aki�E��z<b�<�h���Uƃ~���Y��;��WE_|�����"�3��7t�6��㕞V���!� �(��'��iy,|s��BQ%�
q[}�9�BA�B�ч��,���ao��4�7��UDAEs�}&f�� �}��z��&���r l��\�'��� R��UU���U�H3�O�-��N���������D�k~�³���������9�_A̓:�`?q�0(D>���Ӂ^ Of�_8�I�N�������*�&��|j��oF��z�x`� �T�O2��a�4�a�i��I�$���ͺw<5�(���C�G۝���〧����}�PR}��
kK�s����XsX�q�1M2�� �������Y�5�� h����@+X�9����>�?|:�ED���<j��c&P!�~qb�TߜtS����ծ����l���F�8O� Vh"�x��dřT��䄘r�#G�EJ����3+>E	�
"��"��9��>���=����_��8oi��;� _��+\��@�v�O���RY������d����E�r�P�e�u�9��v�����	A�Z�!ȪY;n�h���S�Y!��w�!����9ϝ�5��I�� �f�$W�Lc�ʳ'�֦�*`x-�ӻH�s%<�l1j�Ґ�E("g�Qo=F�-Q0p��Yy�F{�2��9Z`w�����</X����, ���1K��BbEJ�
@U��n��e��7L����o
P���|B��X2h�/���gǲ�<��1+�?]wt�GG��5o!M� �������k�5��f��0��y�n&M����h̷kw+���QIZ�r!	���+j`��ދ���Q'o&*S��1 8��p◳�Ii/�+
$TT�8%��Ș2�"�Ej���15�����ۧ�gݮX*��k�	,��IV��e���56�qz.byɧ-�nB�Zu���������NC`�a�Z}���b	��N�.��Tv�y�$ZM��.g����,%R$��9��9�B_}\�nш���!3�M�N����G4<�=tZ[:��k[���e��:�klZ�T�""�}@���GO3���x_T/~�?@��[q~f�VV�d����CY`�II��l�l���~�>����X���wW��#���Q�g_f0y�*$}r�ǃz��P�?N�Ѡ, kG�L��2���_1�������)���Nl�G&v�q�!��Wiͥ�F�
�E��� ��#��Ԙ���E�2HU'.S�i�ڃ�w�q����a��E,�Lbep�۷`J�{K�#��=�_���v����VB�M�����g��ħ2���qkoC�o !|���ί���/k R[�/q%��艰�P�g��ȩ/IS��ئ�n`my�U���px�;v��W�8��m7]b��?C��L!|��E�$��s��<Iq(����GL]Ѓ��e�Y]���:W�c��uX-�$a�sCp��bD�ֈܡ���W{U��W��E�FF���:o��o@I�z�0Y�
:�6��^	��Y�����i�H��[8O��v��Ʊ4e�!�Gڌ�����&5�z�굻�^Yͱx ����8M�Z���ˍ�a4NH��^ӡz���ɮ`I�67���Mۇ>�J�\�hN�d��3����b��q��;��?#Frjo�Ӌ5Q>��+�=U��}8�yh%�@BJu$��i�w��H;�|@]�� �t �؛�xΑK#v�Ey�y�jHj��i"`�	��7\���B1���[������������r�	(�f�,h�Cn�Ҽ���я����:�o?It͏zT�%`P�̼3H���Y� ��~�*6�~��U��"r�&/Z~���?��̜�}������0�@�z������j�!�� ��A�i�a��3�ǩ|�$�%g��kJ>������x*s����l�D,��a�g��QBH#�ƙ/>�U�jIǎ�oƥ���G}8��h��-�k'㇒N�����&�!`!���@�6����n��@a� L1c%��kv������:�'���?�1�����7�w�v�)�Z	�]z�;�w�����ϟ����g�B��yUL�dK����e��+�(+�)Vj6�����B|�.�N�7Ut�Hov��B��͐{�w�}��@��ͼ���mԬ������3�O��	��y��69�8P����	�B��(���"�L� o<���_)^�����s��J��E��^[+�QA�*s�_�d���W4�l�"3�Sr��hxMb��-����x��%Y����B���`߹\%s<U�:��xƉ�E�l�z��%�� �Z���
a2�Ԑ���}�8��3e��u��߾c���� ]r^ҝ��r����L������(�06M�zkSNpI�l�#r�o��)�ӯ�I�9M�_��=�AS����z|��f\K��M{��0|�U1���+	>�6�x�~}��u1��Ƥ�bȺD[x8H���FT?z����i�VϢL{b�x��I&�o�^�Uگ���n\?}�H��,Hص�j'�Eb�p�p�B�kE^aV�i�Q�(�8H�\��Hf���*ߢ��H�ͷb�H�v�ĭԈ�xK̓�y ��m�Ċ����}�]�Y����f������+��C�-jhd����Ǧ���`ֺE����o寔�{�〾�H]���M�0q���2(�?+� �@
���y7X	>�^>�z���{�e����>�$����'W7ׁ�8�+��z��2�0��e��Α͌R{�	��ׂ��&'���U�^F�2Z���՚u��' �=˘����Ǟ����e˺&�ټM)t�7�T�@��j�������n`�AXl^�A�f$�h��n�\h�L�m޾��Upy���GT��,���Ca��ګ��eL�b\�N����9���ex��}�����N��b�e�A�����S6���=�:�)��� $;\�H���Jɘ��Ũ���%'�^s7�X�o�?��Sm%��U�g	��c�s?��/C@����ˏ?�qQ��:��&>�w� hn)�&�t�J�+� �H�áć{2.aw���j�������~�K����d��� �u�8��S�Ɣ��7��KF���(r����V��C~#<)atc1�����"����Q偓���^���9<7��\�����;��F�1��h��L�=A��ށ�&��}�H��b�w� =F3�$���׵I3��On[�C���K�~�~�k�?N��`/)m;󇓲�8?��P:j�h2�`=(��H̩��
sڑ���v(�P��U4e�;����BЯl�#� ������c�����ϯ?JR^E,_>�~#�n�0���0n���Iq��.�~ɧ�> �x�7`�c��nwQTY�<�5JE��ͰǷ��H+���ɶ�J�Aq�����܈N���(���5�b{�<B�I�����R�ϙ���� �>��7:d�dp庄��F�Ƽ�9��R'��[��-�Hj�&�]�g�?�5(�4�~=�;��X%~��	�Ɏ��¥	?����bw۪�m;C���ijɆ�$�$ �ռ��js�4���^�K)��M���$G�� ^���xB��E�����,�kۤ:�X�F�?�O�DjE^������%�j6K�=Ar.c>r�P�r�W��I!��J�Kl���GI�@�����y�Br���w�/�g�'6�G����~HY���@��m���>%v��P�_�n��{����ϵu,��;�ә�
|((+Il��g4��"�x�%f�6y���~גcSCfMs����'�|Z�".-�>�tQ��Zlt�G�
u'*��K?�B9�D!��C�t����C���!w��'�=NБh�D�ڏ&9N���;�ԯ�˙�A���A�0 ��o2�%Q�/�M�����Ȧ5Qg�L������ ��ѵ�u;���F��������\�<���Id��?���i�k��=BnA��`��'3lr+���5έ���$
�%X[Жr��\)a�ӻ�'PR%{@�z���f��3	9��J��P�^$�x6������E4���By {P	��ε�&i�5����gU�%�U��|'n��/�#{������P���Ԃ���ڎ�N��^)K���`� �m�	~�,2�v��W�=3�L���i�3�x�km�2"����kA���y��T!��PN�j鷤�<�
)�$�W��F�K���Ay�%�r8ETg�jyN��Xe�vc��!W�vt��[�2��}�D���/��c�ӷ��w��{�7��P�t���Q��3�b<b�;+�{�uM'.;��+��it/N4Eňv��P�JF7+>R��Et䬇�C/������}�a&$O�Qv��Mq�^���J��(��~���WM��<�ƍo<n�d�b���_a�&	�E��x�G����-��Y�D�d�`S�gcZG�_}ڃ�j��u�0��xn��q�m�t�:g����8�4�����7�N��N&ml��0�콺Ly�ه'}B��ر���0j���@T�	q8&.�pi�ȩ'B�f�]���ދ�Nx��VT����3н�'�˔�������D*pA�mm]��E��8�d��|5��[���~Sy��-�F�ˎ�$��1���=��K�x0�H�_���/��T�R��2(��j	YB�8�tOH�3V���B9�v��������g����+��1pH�}:��!�c˒C�?5Ʒ�3�K��"X(ӣD?L��<�{���u8M`E��|(��ծ��2̩ �@�Ѝ1[u��H��t\QJ�R�[�p�̡����,7��79G��X+9�����Ki' �H$�u����蓅���'Z�xs�I��7c�)��X{����cC	uJ4v��G`"ʇ!�]�����z!�b���������@UR���EH{���2y�܌��5HRnd[@�[�C7��N�	�;=yҰ�"� ҎɝL���y�����>c�.�Z�[��]e}.UM� +�xu����+"��Қx_o�	�~K�`X�,y}$\��/�{&,+*�H�X+�����9��__��*Ơ\�؟������"E��Kv@\��jTV޶3�U!sK�;�퀎������)�w��7	U!!?��U�cLa9�$O��vä����̅�{�� ����r�L�Ӑ6(�@u;�ڭ0s"G�B�
Ě;ЈG�Q�Xޙ�&6Ip�����1x�GbH�qA���`�|ۭ~��|�A�y`�y���r����'#�̞n�P(��u�_[��ls�V=9/?ֹ�5yF��ʜMTMq^A���M�c|a�~,R{��k /̒��
�����Ū�L(���E\��[����{�V�'��(�}\��Q��sn4z�F���r,G_B/j!@.R�4�$q��T7�*0���/��٣�_p�Th˚�&�a��ʎmR���~��g�L)����)�I�J�4_��&�{k\��iԏ 4���6��I���4 =�y"y�uA��Tmm�p���o��������5�H���=��'e�9��W��"kmf�� ��ZÏ����|�ĨT܎���͹�Tk��+��.�u�<�	�.�0U[&��«R��N����5>��A �ݽH��'�Ң�bWL��ũO�e~5����۷�`��mo��&y^��f��ˆ�f��J˒� �V�6���+��;��Qki-!z�Q��md��b�p��-�2�j����e][�~��=.�?dc����y�������~��>����W�|��n���BY�'���l��e�N�Wʁ�Be����2�2=�a�Gm�x�{y��8����r�['� �H�=�Ӏ���4��]�!�$�k�lwO7à���l!O�(��p3�$�
]Y�[!՘�5���+O͹1�]z�m��.�P�������\�-d��<�nÓ�.�|�ZH<�OrfU���Pha���揼��������l�]����Iw�ѯ����������YGV2��%�>xL�<�������R::�7�N �B�����U��kgri��(�7̈��zV�&�y~�4�b���W//C۱{�~]�c �Vu� ���`�	���K+��رT�a���S�8W��+�ĳ�G7�ƾ�������aq�3�W
������ h�B��l��0�TF�'Rv���?�4��mex��4R�~�ꗐ����s#$�K�W�t���"S��V��{{���)��Q�Ȇ$�"��� ,^���_��%e}D2Z�:Ο�*�L�H����Tc���L����u�=�M�jH�yH�6u�S侟vƕ8��j�Q�'e	嬰����M���&krgQX�~�/P�"E�������K{���xNb�IH��jR��*���[��4r�H��p%,�ֶ D&	��ٯ�s�鏂��+x���5�؛[��9�2��:DLZޠ��J�%7�rl�m.�ܾи%
�g���z0�[G1�ү	�-�E��k�Ҷ��袹��=�+�f�m�=H�EL
4�8�7 ٚ��}�q_��S�A��%�4�e�M\��,����#�?(nh> �Ȇù��&�e���7�t8�����l�i��io�Z�fc��֭ང�7���?WEb�R�&���DFw�՝��ե���"��K������hP�B2B�ƭ;�h4��������/ٺ���Bb��ϊ��2E"R�h>� ������J�Iy�Nx�U.���o>������3�{�D�!��~uG�Px�-	:�m\�҂!y��bC�	*�R�T��Y��DTԨyRx�.]����� H ��z�u�u��`8��8 �`SƁ!����;������0�t��_�\yvz��,B*W�2+�	O�A�������y����615��XQ��x�5�Ex7&�ǖ�g��a��7ڊ��{����a��^4��uh����@`�U��򄹽?�^�X �pI6l�J3a�Q���i,�����%�{��i����[�&��
By��f�ٌ�ʡ�@C�u�l�f��7]y��#Eȥ�EbV��7�
F~"�6���ZpjY��2�ɭ��.���Q�_{�7�t'��VS.��K\�l����)'�p8�t�:н��X�k��*o���iIw7��.��yA/&2vQ��{�D:E�)N�T��E�ew����M��H������C��Vf��5h�Ώ6:_t������?G}��`A��)'���|��A�܂Ȁ(�o:��M��l��B��[�ڄ�Wx��O��y�o4#k-/����_2x &���4m�Ү��!�]2�׏L���4�M~i
�� �U���R܅��	O� �+������N�<�M1�![~z�l�!�̘H��߯+g�GV1Yہ&m������W#�L�s�v//��X���bu^mg��ڿ?.w4�+�������S�V�l�4�����!f
�9�n��a��i�$���if�i{ͧ��@�J���;��8h��Z�䠠�ǫE�Al@��`mӟ�y5�q��SM��m�QޝL��ݍ I��1=�*@��_�u0�Ȭpq��m;�U��غ�m�Ko���4��aT�gjxJj�)� �ZhW�/ݭl.$���؏̌��MOZ�Xm�k�c �D!�#!�W3�!���k#�Z���@�<mtن�S��i~8�y"T�ۜ�֩�$�����oJ�Ԩ:{J�$�3Ժ��3�)���m?��*m!��y�����E9'����͂�$d���{�1���|R�[@��Ӗi��$[P8�r�48ҀU��&�9qo"AB��rUd�)��)�Ώ΃
�֊W؂Ww�Mŷ��	DSW�݀��!���ceh���ڰ
�)'�{�.D�.J9b�a����[�ݔ#�*��B�ru���4�A� �r�(|kg� �
ɐ�!=�4��P4�q�b��c&�D[��T�>�D~�"�ٰ�4�����e-X(�T�/�,y��%4����r���zf2H��#�m'|`�1��5Ӛ��U��6&e�a�c�$�D=�]��� ��B�_}ƹ|�����_���Y�Y���8K<�0W���b@��� dL�5���5u�P��I�"׿T�/ɭjF�d0'�ܭ��N4*��9�k&�v�5A�:����).��5 �}[�,�WepDI��X��ZS�L,��ۃ5�횾�w=��D�%��'���5�Z����$�_HС�J�;#�|����^*(�52�n�-(��'ٴI�w�z����0T_?%��Ԑ�!2�d9o���P�.=�駌ր��(��e��/[�鑋(�I�6$��GLuy@:?��׌�|��f'S�G��Ι.0������B��~����jsΣT�6�;�W�l��U�ߥ�T��4��88��3���A`i�YLU�A��d*�%����X3�R���J�j��6�[ϫ��m�b�na�(?�l�H���S5���>:�U�\��];��F����Ufъ 8 ���	QD�U k������щ>LC�"��4��Tw������)���w
�6m?8ు;ϻ��>%�TX�T��{��k7n1�~�-1�D�
'��������dK�c}X�mR�J�P]9���D�����,na���-��?��;v�n�}~۱��1�REA�Es!�ҵ?3��!���+���a�;9|�	�����V�L)B,�\�2j'����4B�`n��du xmb�w�\���)銴�$�0E{c3ZodӉdH['�ʴS���c֑W|}��Kg4t}���6������������7�_�0�`���~߾�Y�������cЧ�^�����x\�=��i����pd<��:�^|^�	h��K���4媡V�fDu?ݼ�����V��a�.*�X�����ܰ8:�@���Y������1�bc8:
֠l6e������1���ٝ>�'��N�:�N:v�~��jv�%u�I��F�U�E���v|�a��<��I�/=4�K�6T:��u�z�{��a ����?YZ��$�m<-�?!F���l��$�b�an�F�J�X��&`�@�Rv|���yhv,���sC0�d6#��F�>= ��XyG0*�&t���L/G�I�H̽-��[���e����C����dA�~?S�+|�26w)�q�`~~C��p����oFF�	�
ј��q'f��=ǿͼ���}:���%����1B�ʨ�����I�u�kJ��\�0B?�
,P,Y0���'�Tz7Ȼ?��Cm-2h) QKu��eވa0�b��CP�����,�����P�)�Ec��2����"�yG��}L;������J^��=�G�:�h�F�U͘����h��Uo�p��̵_Hmi<<��������C�ŷ��/Q�8��lK�߾�Z���պ0Eq��%=��/�1�
r
����������
<t��׀���n�X���&$�Om$&��!Qh���Wd���������^
���Y�+9T��+�����}O'y�Q��#��K8���G���kˌ�N�oU��8)��Z`�r�p���b���]�2�����lߡ��[���03U�ȼ�G��V��O �,�G�t8ÿV�;bvN|*�`GZ9?���P1��
�K��d׹���� ����n}�g��4�d��q ����$�co%l���A��␎��2]��ܣd;��P�נ״u.��u��k����?���"��V�O���CSa�.#���K�G/`�<��5w��g��4eDڨ�鹲A�e�e'��̘6���`]-�OV#ú��
���v
�r�`�ҵ3D5b+(ȟx��� ��hn,É��ǧ�[�Ξ�G��y�B��My>g�X���C�2�I��bQ��Jj��`�f�K�x��������@����o��Тy�D1V?#��lMM�`�}1�h�kε�yJ6^Dv��v��4��NR�vg��Hw�45�F�B��"��ٍ/J�<��å��0��z��
}
�h����)8X(����(ܗ��g��js����-�����򉋺\Æ[E�MK[��JTO��+,��^��:����M���q�8�w^Z5,����^�Y�b'Y;�$ަO����5zpQ�*��))z7�EC�Tc� ���� EZ>���.%��@n����X�Z��fdF��U� ���R��4����o�]�m�}�~�H
�����%ll#e�5�p�!���h�@Z���"��G� y5;��pH'Rt
��O�_Wy�f��-�H�Qhs�7��U'�˧����	$��.+2ŔȘr\X��c��Ԛ���R�D&0rm�sN�f�)��ͤ�5�H����(��3ܑ�z;��IK� Տ������ߠ�H�ͻ�z�.�]{5	qdy��Ꝝ��\�a	�^
���0���@M����ˈ"	��$��ir|��_��f��E#w�zq7�M7Tl&W����Ho�~G��ů�1	䬌{TI��`�>)��q��M"`�W"�Uta�ο`>��ȥ������𧻓���������C3�rO��dJ% ڈrG K�+�	�!�������<��"k����ލ�FOi��	�SQgx�u�3��f�V�S�}���~F��%wLgf�һ��JMV6�=*�W�pJ�n$ (�m,���:"$#�GF+R�Y�i6�&�7��2$hT@/}U�'#t�f;�iI��ܿX�v�o��Ou�~;�m�e�;��~�y��@aN�MD���n�{��� �8?�
��e���x�y��<�"�Ws
�!=�� ᷲ_Y�i�^��:ߡ�P�	UGc��$-=Pf�8ck�d�7�n��<�j��y9�s-uI�h���/'p�c�GZ#�i�y�S�Kաm{Ne�����F�̘4s�B�̜R$<�R�Y2�W�V7lVhnE&&�,��h���3�.jY�)�����XD�[S�!kWrMgck���'c`K"I�("4xt/J�Tg��Z��ֲ4Χ�R3A	#��3ͷ���m���SxO������������Z�(1�[�	���M6�(hpa0ܦY�k~�M﭅�!�g��0�a�v+��QQ{�$��ŕǱ��<��R���I��MH��wAXd��끇4#�9t���s��}��4���ɬ�9�G�U'�NgD3����e��%��8�(����� ���H�Y��`x1>�[Ƅ}���0Y�E��CZ��߃1��)�w�>�8�g��h���$/
�U��y�kvE)a{�q����zz�����G=���/0���r�1<p]^�i@"v�^K�X{��0��6�C͕6<����H���`J���I�<��5�|͋:�M��u[� �^r��=��0zq�FA�2ە��;z-;�p�I4bio&X����G?�z�� 3���Q�ʬ�a�C}�24�"�pN�y��29��Y)w8���1}���Ⱥ�y�<W,Qa�;(��t��ޫ($�ú�S�\�@2���a!���r��4���)��/��͏�"Q���M�3Yv���L��B�ҹ���JЭ�ڃ��;�p����.{و]0�w���b�;�$J� y��q�Tv_��Tl�!�pNPְ�!�>�aG}%F2�K���h���#zZY��>Js�x����l�qΕQqh�P�%&{_�Bc�똗ٹb�Qk�4򪂕j/�*p�O)�iN쑏�LR\V��d����LN{w;D=�>�,di�5 �\]�
 �N�&3���q�g[�S���f�ć���4�Ƅ,)�OH���iI�S��$��ϟfvڱީ��bԹ�䁛4 %���N��P���:��0�%β`I��ƅ�\�$���y�ܐ�:ߝ9��Y�e�A`����_�p�baW�Cy�q�� (��r�ؚ��[K>����	�*T/g� [���ׇ�4��ĩ�K�_M�ad�N�Q}ٓ���b�0I c���qib��oN8\1Y�+��"2O��o��Co_������ҵo �X�e;���������	��Rr��sO]��UfJGM�0����}��G��2�V�����:ս����o��:f0���N�]�J�D�Ц\�����ǐ����������:���w4�2�R����&�$m�)�e��|<!�������P�x	Al���[([X���g���%Au�>�O��E��v/}�(*4Ÿ�Ǥ��S�W��4 �*����'C���Tc�'	7�����#��g���)�9֟Èb�U5ݩ4��؛|J���N�IA�� ?^��+�& ��c0�_�k��Óe�`RщȌ���6'���$Z^X�YH���-��b�#�;Ȗ�T"!V'��L�69])WN�*A=�qO#/
u/z!Y���g���|QEh &�V�<����y蠸��e�|����GJO}�_��w؜�KJVP�e�(��|���r�/��������"��_���s5�A�p� 2��x�Z�j1$=�B��,#TC��|�g��+,'�����Q(�����iyKԄ�j�Qp�	Bs<k��v5u��97O�4�5X�N�
Ff;7���ʞ���k��P����H�B5����:3��(�t��7�vs�<�1-�vQ����W=��<��)S��k:/mwi_ �pK��z�L�z�vX,�V��)���훌�� �cr�==�w�D2��+N4�k���&%��㨵��2Ƴ��\ĉ)�%�L���No�N\��'�"�st�J�"$eb�$^�H��6kP�I���@Z8S�)/��\,�'� ��s�wxt��彎�N7Ԝ���CؓI`��K��g�6�5.�����N���)&��FN��P1�sIt��>0v�ȥ��-�~$�dj4"E.JIG=1ia7��nU@A�M���f�����7(�N��)�$f1���icP��s�9���F�Tɦd����5�AA��)Q�rFW���%�ч�x����*I���^���>�� �A�GH[�t_gՍ
<�`��w)�9<���l�^m�9&����7V��b�d�w�$���.��Q��w����!հXVu�#U� :4+�xq��x4p��a�9nm�� ��)��n/l���В \���o�b���9��žE�<�@lfd��&I��WkcbE�F��Ҧ�b�B.	����<{�~N���.:�b��u�p���q���X�+�C8 A��v]��_����[�9��=+���2�3���W�U־�?=��³��$�r�G�]����g�!e ?ܳ�j�p�ӕ�?>�}����J��/�&[-F�pʤ0%��Ԃ�g,`t��w�4E������D9���M|�
JOґ�����"��`V���@�Ϯ�ݟ�a*J�U�H�u&�PS��_/���C���q��1�h�	P?f���/��@<4��j���,���SO����rR��;�=��+@��[�,�ҝl �q��Md�[��YИ�qh��ّ����K1։���0>)Ǒ"UZ5 lF�y�Rm���|1�kAd�J"
({�RP)�|���-b���#��7��$�,ff[`n؏�Yx�41@N�����q�f�A{n�k����m	?}R������z"@����}|qȄ�z~>��������|�U�t��SHXe\��柽�y���@':�2��O^��I��� 1��c3R���W`Ԓ�ה'�i�N��t��^P��Qd'u��DU���V.?�ǡ��ThR��/h�I��ěRh3c��Bp��pS���� ���,�bݼ���:|m9�j��^��͝�.���O�M�O���o��ǣ�w6�ܞu'uo�m���oV8Y9i�W��.��=AF�@n���B�+��u�����A�a�2Ӈɖ�3�qz��L���'u/D�?�R��P�4��pw��dc��#��2˓��1�E�O�3	�7�g�����|�؂���W��4W�z��SEȎDR��Í��y;LϿ4r/4�8
QV�ᱧ��?��L�xj?$�m���^�1�y�Jp!�%�P^��ׯ���q��!y�Y����J'd��tL�\�EH�Ë��5�������{��WG�6��6�����ILIN�R����`oʢ\��m�(���[����~P���&��[m7*��Zj�]�$c��#�����G�2�w��l|���y�)�����s�M��--	��}�+îβ֓VNd��5ba�eK_�4�@�+ T��ퟆ3��m��?zG	�8�]�CjFl���-lܰRt�0~69������'������	#��3g�z٭�U��႗�h�Ƒ�� �8Wu(<�K��!�¶���]��7�̵�U��LFg�_5pt���J�1k��(cl����-W�5�ޓ�X��D��?���+�tc.SRjAe�	�C(����*���9b�M[�3�0�(h�L3�%��"�_z|\�`EM��bH� �o��%�NO����i�`�5T�\o�)�%��{�����{a{���o�����F��DV~q��-{�ޮ��T,^ysH?Q0I�D�1�sG�T��<k����.�3�A��r��h��?�3bnE��_<�l� �1���qp�lj�%�<H�SҠ�Q�g����dKfjq�X�&U�ن:)�>��I�tI'��&�Y�\���}T "�����]�N�M<Z��U�[πbi��%���-�ԏv��K� O��x�,:��23���^"�$ӓ�Hp��̈�0�n��f�:� 9<�55�L�c��ҙ�y�$7J<����4�����&KL�on,hsZ硿żw�����H?`�$�gc{��u�'�L�r=}Kĭ�6ԳT\&�٨�P�`�{������"����N�<�E���!1?���4�m���V�ۙ��|Sߪtd�y��H�v]l��H��Vl����0]��7�հ�^aqD���'s�2[k�����w�EI��%��P�gU��}#�\P1� .�6
8����ԇ�'}�kKG���2����
�6"_Ⱥ��z+��k���Cļ�_�陋鋑��+�w��@�R��w��@F _y��f	��qa-���xL��HD�|�Q'����[�	�@�X$1Cl��e�6;aX�Y��z��f2A��]p�]��7R=�O1���*ޭ<����އ�rN`e�W�R�_��ɠN�A�B1G��)�6c�>�j�z�}Ɛ����nk{��,��	Ӭ��Lj ��c/V����p�KӰ����7�pEL)ܔ�x���H��T!�m��ږ:�(�?3���T��k1��ԋHy]H���#2�
��-Їw�4�]�'Wla�}r�yB]�̛{�E���L��^V�كE�9Λ����CׄȮ�=��¥�"
����Eŏn��~��h�`	,ΠܷeS����Å�0vO6�_��'��L���F�D��^�5� ������غs�/xq���jǦ���ES^W� R��U��`/a�(/��Ϯ^͈b���&⸫$/�0w�Bw���e�."WM�54���9�)���q�R�ǖf��}��l� TCG�+R�5b���O�9km�n�嗀zc�����(>YK��O�4��@}���M<����ؾ7��<%���B\���s�?M��m�N��f��qG�!h��½�|��T��к�}�n$`�z�l$��&��E-:��T�P��-�{����ߋ�au��*�-!���D`��#D|� ,F'�;A=@�N.�IZ�����꼬eԩ� ��]�SС�,<B2�s�O{���Dߵ���O^B�}ai6k7���Km�o�gc|���96�߾�U-O�A�b�F*=aqu��p�$��UAl������e ���[�Ԉ�y���2�$�$���r-���&T����l����A\��̶Qj�@�_���ԤMfKW1��Z���/��y{���/b�e�?R�����e�n�U_�RAwm�Du��O���ah��y���!T���3w�'ac��A��r��-�U^��u�Mf/��HE�uHB�E�~�9����Tݶ0O����H ��\]u��U=e������>ȉ���bl�W�m�OǴC��bH��c5��_����=O�􊐧�E��1:�X�R<`��+�*5�IY<�0�7jF�]\FA�\����Mx3��@�	��!z'���o���\P	龖՚"�������ۺ�(G-���	�-(@fvX�FZ�h���f@�"o*[8A��#��)':�ߧ ��<c���]aԶ}�Wb.=O��1�'�Oq<)���m�2��'������X����[Q׆�׼����dj	>z� y:��ୈ��*k�e������7 �e�Ʒ���.���OU߽�8�z��PwI��G�w� CFԻ��N��	(?z�E��t���F\/|;F��  F#��� ��,Ǫ!H⺦�ǻEʟ��P�-��+���7y�	f� �@
J�ֳ�i]�p�ʹQ��U��7����d���=���fl��O��I5�Q��zh�
�[ޫ��! �<bԑ�A���aJ�Ă�f�z�*2Q���^���,7�w0���2��s`�ݰ6:���"	�u�z�.Z�5\[FM8�eѤ�{��j�T�N(?_�j��*�2S��M�I���<�	/�Ƙ�h���D!+�fz��.JA��<x����&�DմI�ط#ΩH�1!AW���cO�g�,'a^�'�(�N8��/B`���<jp��i:��o1�<��F��81��+�g��o�����Xn�EZ<b��*}s)����l�,�`�#�ۓ���c�	<�ԁ��v���-�� r�'�/��ȡ����K瓃C�`�vdᑵmۿi�}�r�c�j1=�;lz�[ja	����}�3"��7 ~��"�J{▌�/�v����/��m8ޱ}�kЧ�����m�؟F��A/I�����U�ڢϴ���H7�TF��(�[A��]�l��fS��5�����ǋ�84Uu��w�c���G?[�3h)S��ktL��Y4�M�c5���N��`�Oۗ�0*@H��KT2�)\��j�P���Uю�����fKV_�����n�m�W���4�D���0������(���a4���E���gܻE��K�����|)��ZL��29��3'U<bhϓIcK�'�h
^L�.�>А��O!�I�)G��f���� �<�3���xL�4]��z�蟦>�����=׺���r�<	�7;����B�Ԣ�{c�H@��r��Z��7�Ϋ�͙��	�v��fAU(��4(��
��G��8iN.#!�%�-�D3=�Q�TD,#�ύi����+���q���6�m|�����(�a+���P��k��u��mr��$�,^��{�X�����V�ؤ����Of��>R���9s���hM�ড়k��Cm��CU�i�T��1Zb�UȍM�s[��=�=R�]��LP"�<�Qu3�(����mҪ4{:5����NU�	h%�^Q[Xgȶ�f�]���#�-����(���u#�<~/�Y�o�82h��Q&���N�6��nn���7ܨ�;d��r��|�`��rq�֬)M�I�(^����N�.F򈲠��~4�� �ǯ�.�"�7C��R�`��!�� ��H�x�(�涢��˕Xeuh�p0�o��3*ـ��.�E>شOr,�)�k�C� �0�h
�������a�P��)NڸI]��b7ξ���7(�T�}�=�M9���L���e�yIe�*>R��l�b��*����FN��n�Ĥ�c��b���$N�e�çc@G�A��;z�˽6v��2�z��]��\/��U���ٔ/fA�.Rp��aB(��#,�|�/o٢(`���"��v.{����R�?�AP9`�X���ʿ�>A^Ĳ���]FHc�z��!C�o׺?�R���8ϟݛ��P��k�	m����mw�JM�9ߢ���0�Q�e�^	+̮<��w��	80���%E�>l�3�����&��Jxo�ep��OU"|
�m\����-D�����	Ǝ�f�F���M�_5�/AL�����/���jXP"w?{�<<M�g8id�,{o�S�e*����ՠ�}C�8��{���
3�2fѼ{"yG���1�%���Q�jO��G9ǺPA���3����6C]��B��#-&"��D+n3p���h��*�m]�$TJ�+&�1(��77e��-��C�r+I@�2�/�ɍ��Q4�ۛ�ȼ�������ϛ�)���R��b�A
p��W6�n������e������F��l[�B��<��.y'w ��4&�Rg�KƧ2�Q�S"֚I�(��W��z�  &b8KU1��_��p��	�A���(+�tX��Jp�¡/ v��4y݂��0+��>�����
<k˸->S�>�&n
 y�lZ��f6����z7Lum��� d���h��-��� �)�+s�ߣ��?�Dh1LqYα.��m@����؋͇���u*.���B}�*[q���_�I�Pʂ��Ƅf`]�Ѩ�
S	,���'6�vN2>{��U�Y敼5K�Yc.[B���L	ǌ���z�h/��(�!�Q�e,'я�]lǋ�:z3��
�w<1 �P�q����7�#��QxE������U������7���Y[*m=ir({fW���)`��p�P
�۠OtcHw_7r�ݼ���d{C�|Ao��7[*Q����Ѯ��q��7q4�{��������*g�QeV��L�CϹݭ�WҦ��L�ZA�Uۉoԗ9�r����}�H���W�-�΅��LAY����$z��jY�q�G,�{f"��q��j7e~�2�
�K AB�T�F̀�����/FؙNcG�j|�ҁ!X!\C	[ؖ�
��M�Z�Gs�q����K�Q�0B)����f����ۍ�s8��W^���#q�����^D�P��4�e�c�'�1HA�z|#lXU
K�Z�*�q�kqbOh�eR呓t,N����� CWe��F�"o�g��
����陮
,A��25�FV�y�����<3�J�n�T{N�Ra�r��q�ޕ�zf��+e)�	s��|v*���[}��0��~��oc*�jC�b�sqQ2�%d�
�JQ],�G!�s/�e]���A�8���9t$VL�C��4<��e,���'�ӕ�X�h[��#i�׺"E�+�1r[�F��kf}H�?���WjP�f/����3I�3W��NC���������1�D!e�G	��ft�܅����&t.մ��I�->�洉��}J��`��}@�����Y%öh}��KG���Ý����|�f�+WD�{c������=����FL!�ٮ3k'�1Ԃx�xc}�!��� �����x׻�F��[�L��!����B�}@�B�N�$�<���z�#��4�N���ۙ�G_�3�&L�� I(]����]VZ�������vZWFb����܅��U�x_�&oy6��ԗ2���U����K~��1�ccд�D��!���6����qG�doβJ�$� �R�>kBЉ	fh|@��M�� a�?b�_�A�5���d�;�&��q~�˓�8HD��ؗ���Z�C!�������ʙ,D��J���';N��r�	�������i��1�Zþ�ޒ�w)�a@x�`Ȍ���<�'c�,�h;Dg�d�$���'�yZ�a^/fi��&��FDf�T���&]�xk��z���ņ�?�YVí��U��8�p����ADq�s�m���Dg��w�5x@u�)���1���P��c�o_$�,��|=��sn�Z�����A�RF���� '&IT�J���Y/��l�*N�6�)6�����.�*Q^.�o%�N���͐�L>��+�����R?-�^k�#��\��ze�
Q�� d(��M0X}Ǹ�e��)Y��o�z�#�n��ˉ��d�#�K�(v�Z��n�Y�y#��ZU�Y�k��j|of�w�zKz%A@D,�QV� ę�]���;BV�I�Y��G-�s=�E��3{>b�����{��hQ"��aO$�o�_��Y&߸��r��Q�����J
�ސ�iW���J��3��\��ءp�D<�f`
0�����/J���%Z�pRh�]��f��H!c[Ч�|���{�\��Խ��Kѫw�o�3���$g+���e����\3�N5�[|��t���O-H�)��y\�C��.o���D�{�X8z+�x��jj|�� SK:���?�_rۺ�
��+��<)�q�ٕɼW�i��ŝ���8��8��cϕ�6	�0�E��:�kpj=�ͧn����z��w4(�vj����~�.�s
����>f�����]
fx������K��
;
�����,��ƴ@q<��Ǝ����f���������r�F�Td�l��J�'�m71_
�p �e���<5�_�adI?[ �u�C�Z0}�h�<����֑z��AǭW�N��u$[�
�UQolu��j*�t�A�౱�ʊ��Fѱ�f�n B�~�?;��(?�ew�{%c<:g�k�k̅��uYlOֲ,��7k��Fֱ[ޕ��z��v������~�2��q`�Y��L�軬�M��D�W1��pwT��R4�~�!��������<�Cx!����#NC��F~3�����ך����g�w�b���:�����se�W�����L��[�ז�ģ����ln�5U'�"�諈�$:ҹ�I�(�&I�n�<Q��9�>���R��5-�-�P 17�2��ûX�����I �*G�˛�E0n��e�F�F�-���~�c���\m	{ХV�w��y��-]�+�]�!g�fq1�(V	~��h�����F�M���J�orF�KIH���.ˏ�$����R�Jo����1�e�E}��I+< t,�@�� i���i�m��}����\�d��m�˽i9�TD��,X�m�Y���{/,Di_�z5�z%W{��1���`ƒ�4�3������>7�e:�I��E�D���/��@j�`�0�c���S����N�h�n�^�r�b�Xͥ�����=a�,^b�X�� ��)�t�L�|oZ��cB���ތ4x�Ǘ�vʄ* BVƖ�EH���S3$��f;[OL�q��������|\�������r��9�Q �o*sh�t���vQ!XZF�V��=�ش�gUO�]��?Y�8j��Wu��p��È���\��n�fV���e���;��Jժ!��0��f�4q��l�Cgi�O��N� ��D�5� _~�U��8zf�&�^�c���B�Abx0���Q�}f��@t2;o4b�a1ػ�5}ѥt��/>���0c�S�ǨǠ&�O3Uf�\13�tI:����F0%��<ݎķ���.�i�$�	z�*�{<�s�Z-Q�X|���a���' �ҿ�������,]���GQ�Ś�-$h�i���I��tV�,��2���V�Qf	-�^�*�9��LFa�3��wG�E�e]���cQ��i�<����D��X�����Ȍg���C������Y1�� Ԗ�L��Tݮ����*i�AC����*�&�f2���a�i��*���7�FZ��Z �R�#���-��L/A��^J�`A�m��8�v�[1.x[�˜@�QLJw!��Y�8��_���ʆC��� �ʧ|���pઓ�#�z8���
��������c��v�@b�n&�S?o��0-��4ͭ����=�f�CZ��R�'/z=7�6��;j���6$4!gC_�=���������|�ߤ(Ir$c�.�ȃ����T*/8yM2��u=�`p@Թ�Sa8J<�9y*���XH߰���C�]\֯�5�%�B�d�;O�
!�EKX1���ȩ�X�(��S���]�Z���l����L���me8�M0-���"��.�������e���Wk�E;�su�{G�Vm���l�AV���#���ZKQS+���]:=��e�lK7��S"�03��>,W�E����\5��:���B=	o��H���/AI�׵��;�d:�J��Z�ۍ�n���7��1<�p�I����o�3^�@��\���m� X�|��7�G
�Rߊ�`����a��^�5��C \���y�3��hl�YZ�I�s������ι`�f���+6���1&udE�3�نsO�����(Ǵ�J��&�%�(`#���1�޺U�7�ԍ��H*�J�}褬������vkk�xTE����;�P��|�����}�''/j���\�Ӧ��~n�
��|��d�ի�o�ɀ39�P��9��W�F�	��W����3��[蘟��~s����:ʌu'_J�'�Gf�$�����sI,��&��9���p�N[�4 j��T��t��t�T�l+@{�Dv�1_h�ld����A ��Q�=\��^�VYн[dH��y.%� �4�C��B߾pUP��G��O�����99Z,�wZ=[!�}ȋƎ�h�1��R��s���,3j��/�sᜡQ�Ѧʱ��Y��,1ҭ��_c0����ɫ�8��a8BW��Mk���8����')���Y�y;ݪ �3붔�	��v��ldO�!��������N�Ҩr-���,�rI�9�;�FeE_�l	�J]��Ohov9̡Y�7P;I9��Ø2�T�>���s#ʗ�1��ѕ�x�,��9�K��JSnX'ڧ��@\��ț�������g�HbQ����}�4�Dt@/��n�	���@�����V�����6x T��a#�B�;�X^�?R�X�7�5f�\Bx�Ws��^9@�9�ؗ�2�.��z�;�����-O��n�kb+ס ��s�R'yZ+�m�p�?��PUOVS;`������T�P�x��EjG����@���]g�!�r�e�ճ���b$&q4Z����sed��?��u��/�D�<��X��6_�4�(rw�;�]����RƜ"D�e��mA�0M��x���:���v���r������'m�-�}C]�r8��"�i /�⻌���־�N�V�8�ax�¾8Ӿ-��({�h"kH�z'�K���{���#d�4�}�r���o��%M�޼��gw<=tvt�����lY�(��ԟ�����q['��=k���o�'IxnOؼ1}�E��&:d��SD�Z��.�XYk�N�}sB���r�N�V�$�{��/��	L���t�q��7�O�9wqO����ĵ�xIb��1��FC�}b]��H�"!{�D�������$m<+���R4>�?K�;*����#���u�ۀ!�?Hͥ�ȝT@��,�Srg�����#af$������h�\V�:��S��pCw��|N(R�������aQd2ҔhV�=�Q�YC#o���D��ͨ~^ʫ�<g{��S����;�������XK�~�#̍�jQ�煼`ӑz�\�}ܸM�[��(��z��Y��xrhI�}�el3��rR���~�����������H_�\���2����6��bCotH*1��1�K�}gѵ����;bԌ.��}�� ߸e��Ne�eR4N>!�+믐.�\��0���Lf�E���:0rB|����ٛ�2t񠊹�)'��p�^-Z��F#RvGSa��K�*g�5ty�t΂HAL���u�N��W|��>��{E_����븫z�&*X��#%�����1*)٪�rN�JȱD% h;gD��ט4״�K��94������ymu7�c���>���BC�4P�!N,�wn��Í��W�{��r����ٮҲ�w���T�Y�A�F5�b�����\����r7�Ĥ�47���3u�~k�d���]7T��ŀ����w���N�a�t���u�J�ꔾi�k�7J!0D��y��;B��=z�crM�~e}��Sg:F�T#�P� yoP����&\��j�C��4��^���60?���)͟��;̖h��3�������c��S/�y.��Cj��F2�3p ��W����?�Jg/s]��{�Y��k�n#`��R�E�W��߹��J`:Kً��s�aC7T�hD�FG���S���m��z��¯�禙��V�~��I�ɺ�����]q{-��W�]3�ut^�j�n*g�_����ٱ��$���qyw���kj9��J��<~��k�m�.���_ˀ%@�[�NMVګ��L�nKq�1:[7Y\��*/Y���Td$`XAyM�ɷяn�,��0sR=�9�&yþ�mG�ȠI�*���d�kŎ�����&l"�d�}e��k47���&�\�׍���S;ʈ@g� �P6��%�^�1{ofg���B�Ge�&7p�Uh�!����%�R|��c��8����ʬ!���Pf�%���>���v��6~{�H�V�t����CA]�b5�Zn���u#�R�Hi��'�yn(� � �R�(`�1����a+�D����������\Q��*^#h�Z�GF[��.n�t ��"�V*�5'2ۡ)����.�Cn?kG��/L���i�.�}89�.i6[q��@$y=;|F�e����;�8���K]:�b���g`c3�}d������=P��\.˓%���	�&��c�D��5����G�G� v�f)�	Ȝ�
�1����%c�X�̇4q6=�����toCr�C%
O���7��K�HUPp����&o�%E���և�/�Lu܎�_z�;X�5�/}9G[�>����5���E\�[4��_:z�@��`�(/�߹���m���YR�\��/>^ �
oe��C�[ٞ����"��Av������Tҷ��1���3vh7h�E�?�����;���� ث��ȆV��p)ՀW\�LB'�������i`b�\ޖL��`s��<�oWF-�\��,&;l%0�Sвɪ�rt�E۫)�����[��72��&��&�c8�l��!禎B���-j$�xս[�x�y�e�s#����.�`�3�t�����E$�Ω�V�ޔ�UiY�	!	���S`��!bv��Q��h4��WwD� z\��J�����/)�6�׹9���`2�"�ΧK����u]%Kv�e@�k�>������5�e�G�-�ũ�6"��(�Oɜ�)��7��On�ٹ90w�/x#ZD�_�,��􄾵FIXkL��$�c����b��&����@�֔ś�ME��K��	�r��n�{�m�y<pײd<���n�6��M@�K�l�i2�#2�|��@N�$��m����~u7o;Ą��lki|�N\Z-�?b�% ��hӯ//�.�}?>�&_� ɖ��yC)
��~a�y�S�B�}�RA��~�3��J���y�m���/ߖd�������Bo`&tdbeP�����Zi/�Bm�ǥ���K�U$��ԣBmD��O��,���8�EM�|�^T��S��ho�D@\e�v��)��� i�v�3��j�|y �L^��~��,��?n�ء-c2�!½�]�R=/��n4���L�O�2��>�B���)F�{ܽ�1�iRC}JV����H���K`��q���L��)�v� �6a'+�}
^]�'���gKtfr�ZO�K5�$�l�P�AX���S�_doьi^��b8�]�r><�~(Xw��ԟn���
��^svcΎ�n�u���8���}�������&�n�.����|A�І����������,W
N�������sVX��{W�$�Z��t�Oo�f�̲MU���T���C؜�}������Q������~�FQU�� m��C����S1>Y������������[����c��GZ� ��qL����Ԧ��T�x��?��WzkV+B����/���}��N��XO�U��;2�D|�E�u�\��߄�C�ͬA�p�H�d�c<������ph��UO�w8W�,�;=ղ�0[��R��j�!�e�׫LS���|Y�7B+�^2�: �0l�N#�F���C��7��qߡf�2��M���pI�3�Q��\��Ӎ�`�Ԥ�%t�h�Ѯ�P�����7S�����xI0��~S����"�iV�Ĳ�BN�{�W�ؒγ���Ac<�	�l��p�M�NP&4���A��C�}��W�m��a��๲��)��Zʜ6p!`PQZ.�[����\o�;!��Ŀ�m��v��g����'6X8�;D���s��i�0�|9�������T��\��8�Z?�Q@3��}��bB9|����vU���m��c
dR�]갍Z�	�������O�]�C���ҙa7  7��0mn�B�7�!��4NgXx�2���_�?���d����KE��]S,�4�.�H#݉�8�v\$��X������O����Vos���kY��R@�ܿl'�	Է�/}"4���6���ȌO5k�3>�u��p�8�Ri�{$��"F���� �70�Mh�mm���"���J?�!de���!�ij�������e1��6�C#���}����8c�
M�Pw`�ឩ��P�Jׯ�ϝSqI��⠇�X��H��xX-k���=yRK�U��١�a)���}Kʉ���P��&2�5���7����\$n��H��[dj�i,N���
�}{�B���~uŤ����$�7_�]���_ƿ}�3��r5�9�SY��+w���S�S<��dD��K���	
��p��P�'�t1��tC��s:�p-탚[2W%m7ΐW�Eh�l��/ҏ��y��.��c�@��Oy���Ô��kM�F�'}ߢoXc3����eSl�{0%�� 7�a��珕
'?��8��N�h�'8Bۈ�rs�^���"����-w�?ǾM-ul���r��ᗦ%����\O':��~�$���c)��!�������~7����6��i�e��W�/}�}%�RU㬝 �@����i���n��O � �W��(�Us\�p��ϩ���ɭ�I������0�H�ERN+�:�����e�u2�~<�b��O�J�r�-�<�>�6�`�P��u�-�A狘��S���P��"��]nt�ț7v�a�\�W*(H|�`cC%�I����j��ʿ��7�>F
�b���{c2ƪt���郜D�2C8Qwx }���d+h��>hǑ��8���;P=�-�)%�S��\ 21�v� �N��QpO^��p��5D����V7̈�nqU��q5\Hc�_��e�un�*�&�i��g~�P�����A�!�`�q�Y�_6��Ʃ�{� ]=>x�
�V��n��0��ٰE��(4x�Q"��f=~ӊ O���4����>�v����G�$ĥ429Ż5r�c�*�"|W��7uFuvT�ˍ����)yxB;�� �f�\�VA�Uk��2/v?8{�?6�6�S��O��/��[��
y��J�Oj}�� -5�D&�����i�[��������+T�����h6���p�,zKc�}���E,��b;��.m�Q(\���ڐ4lD�*P� �W�˰��m���|�I��"�{ݓ�������q~�����9�:�t��l?4����f��*$��L31��7vr��OZJ�7��"����4�Z+pH�dPj�8 r\8� ��,�,�Vۆ<L0T�8�"��������O<�rl^5����~9�ۗ��2�� �����e�UN�*'�����V蠭w(�kF����]$D� �ٯS-���f$-�7{18[:����)��֑����_�0p}��-�����6��;����O�Ps�`0�g�|zo.1�VN%�0tqB��ㅮ%bj>�?iUb�����a�z�{h@m�洆�q`��nE�a�,��¼�Ù�$�o�!����"���>�f�k}i��4���C+?lXIS�5J"}[�8���}S%�Ύ2=�#p	�yV����Ye��u�n,L�N�Qb�3�^Ԉ��YB��p��"�x_�4V�bږ!Ri-O�X��ќ�aT����;��2f��2�����K\�����@�#�������}�׳@	���fAGI���kl$�|�NH���'l�P %����H�j�}�B�U�ѣ ��e��Q���zC��L�s�{vt/˹	��}z��<��<�f���[�25���k6i������`Hhv�'X��H[?S�����L�/Dzq/@���hUMܡ��^( �N�յF&R�w̎W����TR잌�V��r�s��A_�/jאH�!����VG3�ɦ�Q�h��GaW�'���:��O�c�y�w��qFN^~,���y��v0�@?-�[Z=�!����W���.�X��:JѮ��M���m{�}:��f�Yq��bq.b��C�h��ƥ�cд���0SW@�c:r���?c� Ɩ�9�y�&U[˓;�,��;2R+���Z�q%3&�'47¯�8Q7�˵��k�Z�Ѣ.cy�0Da[= p[��L�Cg��et�7<A;�M��vGd�|w�'d,�Ip�i�H�A�1�N���$�+f��[�UlײXjZk>C�źn����Nl�ן�P�G)IC�;y�9z9�vͱ�g��i&L?��:�' 1�3p�ӕ�ht�!��O����Z}��f��|8�;��Ud�[L;.\�N>��l��I���=s�O�G�����@sm�pH)e�5h��0��L�`_����r�t�&Jcͱ~i�~��]����@��E*�ըk�m~FŚwg�p�I+=%Hu@��ث������I�����N��������#��
!�'}�Þ|YI�M�bkc/�'zwNp����[�-i����{8�(������R�
 �O\�SJa�:2���Q�+O�;�p&�%e����xv�!@r�Rآn����>�����k�c���À���}{g{5�Fhϕ�~yz1�X�¢��4-nY�8�#��],�gr7��J��[n�8WN�u+$4�;�܎��<ܞ|�!������ĀΞ�Kt��[ʹq��������֚�tONj��bvN��)�Hмd˻^�)����S��*�.�������_�>�j�e��[K�h�c��:�xu�3)}�w�J��>0�D�DFıJ��Z�%W[x��,������%�;f�����3���~��N���.�JW?��b��Q��`�e�%�*�Pj�$d��_�&�_�`�؇]�2�H_<-�$��o{����Է��x�P��hi	c��~`��W�K`g��/wֻnlj�>��4�[:�=θF�\���/A�,J������3�e��I������b[�Z��/�ۨ�a��][CY��d%�D^aD���o��k���t,1�u)˿cl��m*��U�Yt�~�J�%HWcR@
�F���ew(2T��7X��UD%>�)�e-�\禢W��h7g�0'g0p���"+����'�u�0��#���u|am��~��3����A���i~�D��e:�NXq�=*������;5L�{9�T��u��}��륳�&��2^��:��+�����v;�Ā� ���� �f��bginO	�q8��^����y�V��rB�����h8���tyd�"2HC�t�ǋn~M���2���g���u�_�o851\ǺgQU���M��E��!�������+����2��<x.�_���53����c̐.�)຤6����@!��h�sPm�#���W0|]H����kގ��)���>�De�����7��T��(�x����wX��=La����qgs�nx�դ�5�w�N3$�*4�i������`եQ ���mmfYE�L"�y���
��^�:n��&=��`�۞���`A��M�R=f���(霈��0�H��-�%q��Ӊ���1�;�]��U4�����S��	|����ߨ}��|ק����W!`}�C��dak[��f ��$��-��\N5� ����l�侢�YК��,���-�rlq�Yb�
ʀ^m6�Cʿ�G"b�Ꟈ�1�I.��vLE{U�<�۞�I&m�g1I�?6k۟V&���%p���������<�BIr�;6sx0�r
�o5m��MS�h�^��$�%˦F�W�e����SI#X;q4�eiu���ڈJ_��,��- ~z*�;K��9�7�Јv�!>Ƙ��D'�H�e���:6�y|��0� x6(�vp|w��R�p�';��\m{�\�TE%W�h|x��jţ`$\iL�4�T>k':L��F��F�b��]Ԕ�����>\Q#55���?J��r�`�O]
�ݓj�o~ ������}H�����Z?{�a`Iq��eǉ�}#�[^̅��]�]O�e0����{B�
r�ߧ�C��W�K���9�E�+7�N�&���h�/7ұ��kj�
o,���� Mi��~7N�����7�B)y�?|?~��[��n�	�n?Th�5ob�~7��t��O3�Lvrm	~�M�����8�bHy�w�d�Z�0]�w�������Ĭ�+/c8���J���:�<I��w2��1ecf�v� ��;n���of��MYkv��]��
wm��t}{b`���&�D�����ݛ�tC��1�e���t��t����FvK�+z=�t|ÿ�����!��>�I�,�_dTF�g��X��#�I*�U�]�xF��k�9_�o|�So���RGi�t{壠D?�Epo5^1�nY����@H��Bmo�i��Č��l?M�oݐ���w�L��-̇��K:ѯM\	o�kQ��/vzHFR�n�,'Z�.�t*�r+�����/�'�"G�J�}cpR@vsB��[�
�v��b�a=�^:s}a��@ӛa��8kr�Ek��G�E;�8���RIj����K�i�ҰC���K0�}B��Fe6��w>��e�M���{��Y���l������9u-�0�ΉM֝��x��R����ƙ�xw����B���7��8K��AR�AW�i+Ν�-凤6��<����8ӕu�`+"�t-��p&�\Op��D�|�3�&!q��ʱU$Wu��Ɲ����Y�����Q/�
�]X�Ȭ��%g�DV���M�vqG�g�}���%���k��_�"ͻ��qqZڑt��tQ�*�Kͳf�@?yy$��:S8����P��"��d�(rB��2U�R_�.�ֽ��|h�5�1H�;���Fk�?X���Z�?�����퓣�c�;��Z�U�!�D����He��Ί����!��D���g��^
�˯[����ݜ�ɕ�ƺd��\ޫ�,�V��سr�M�h@����G�����7��J�^4�l�����0ߔ�W���	~��'�iֳD7��P����u"1�[9/G?�z���m &[�!e�'�6��U����y���V�q��-�c��L94Dbv#���EY�p샸\Y:aS�u���Ǵ8V�F�G4	46�>\�˴���� �[�bJNMO�=�%�#Ҿ��eeay�!��m�K�Վ���i4�ƅm��/'XY�'MX8�(3�׏6cS���ݧcՒ�'�`���&J_;��V�i�2�|.i��_RF��m�� M>����{7#8y�.ś�:��2��5h�Cʤ�O�_M�[���dΤ��!����\�*�x�,��5�UuߥkQ�N���r�b�Ӓ�4;M��,$�{�9*����a���V�i�@"�ؚ5�yw������j��i�>a"��;��Z�+��cwR��.{so����jФf}��4r�sŧ!B=$}�f:�Uj����Ǯ'kq\æD�dԜ��,�TI��ieЮ�h3��kzxT*}����9�mC���l��<y?G�&Բ[�t)![��)�a6LsV>��2B�w������n��2�-���r�Q��Z�>-pk!�Y �΁�q �.
���ތ��5�x	�&�8���	˒��#\@����{�:#�!�C�؅�;e�I��,�?�7I�~�� �*<��^J\ה�܎�����gL����$K9�#$S���Y����F��袹Eh�I�z��}�v�A�l���K���N�Z$Jư�ր�/1�9�T���r޸�ĶwQմ6�-[�����ȥJ�Ш �=I��X��m��"�0���������+�ʺ�I�kM�~˓��R.�'-M�"�EY�8�T\שu�䂾�F[�� �ծ�\T���`����j(�Ȱ!�O��0� ���<�U����7���������=)F�I]�٢j�9�()���4t������x���o$U�g�so��f��������~[[HE�13;;T2l��o ���Q�`ơ�6�L�6���2sm����"����~>���YYPK�D��\�`� 7�%�E��Vt��0=�>)���Ɩ=�ْؼ}��z������m�HE�� Oa{�)�j���T��3��>^E���E�0��Qhɒ��@� �u�b�v�lg��*�]?�l`�Vv���.����w90���r�p~Y�]q��`���V�5�	�B��A��"���:f��b`��I
�>�ō��������_$�h�*4?m�M������
�j͹�Go����P��ѫ��鄝\��M�a#?���骓hš�.W��0��G����s�fΐ�6BV���Ŭ � �SΓ�v�-�\<7��g,8�}gJjéX�n6+Ւ�xݦ���m&�r�?\Qe��d3�X益os�#0�w�8�����LV-ѩ���k�|奝�Gr�u��A��(#��R���.4�(rh���&��L,`�Ծ
�W�g�h����r��>oҰ�W�������{dSO,�ť�]Z�@��o��k�����P�'�
	��羨[w�N}M�;cHiػy�v!A����3�6؟�o�M�?���� 6�+M-U,��`4����"�~�b�.��m54���o�jQ�K�5�A ¢8����������?�/�SNX(�EΟ^��;}�϶|�TΩ��:�b��R�`	[F�,��X����12lmP�q�0ش� �3L��@u��� Y��*)�-0\]pk�8_@ūm -�NbO|�t�3���!���uܶE*��Y��:,�I����-_l'%����ˈ�"T@8�U�܉O�ΐ٫��þka4٘��e��')�}����ʵ�&t*7Ϟ��!��S�w܈ET��	��N��ɋ��o�kO��|����m����?����G�"��r���X�U@>��t۝kd�I�_Q�� ��"�0���ٳ������[W�.��y�����\�nEbX'J$��q��Y�<�}>�Q4�
|omi`�Ǌv����U�� f-��E���vi2�-g�@`I�o2�ל&���n�qH��������],�q�h�ƍ�i��O��C^Zxb�br�z���a;�ת(����O]py�2'��E�� �Ɩؗ�-j�h!�o�μ34�6�HLO}ĞEOm�{3���A0:JD����͹�en��1'Y~^e.� �����ԟ��,�����6��n�bć3o��]`�;=�~�j�g-L���;��XY���ɰ��Y�B��/y�
�eg{� �mq��m�Y��Q�G�	�'��;	���AI�����Mp�����p������(HqZ�<�ҡ�T!�ȯ���l���M� �&C�_�%z�aCs�]��\\�z��ݟ�4z��?0������q-�LH'�>՞��N㥉K�B��i1]�8����{�c�{��+Ǵ?�輩Q2v�5�Y\x#�j`f\�̦L���<�v��Q���=}	�d�C{��������[u�k��!��W��Ge���[Z&�<?W��Z���Ȫ�8���萁7�$�p�ڴ����6��|�L*9�!�=������8N�=	G�o���� Iػz�].�	��'�c@)������^;J�#�1����X�G-����ĝ<��Ss�`�u)���̼�c~<�`AE�wZ�њ��3B�M������l����8�/���{6v"��c���UI	%\�68�g�����/N��jܹ�o6N��`�;� ����]E�K(�j >�9$���HX�Î���C#�D��7�#`&�Ϟ�b7�"�G>����WVv�U���w�L2�΀b�o�x�����:�(����~����*�D΢�������}���OK;����$��!;�#�}|����)��>�F�N����gjy~d.�b��|P߱1�D�
��C����74��X�$c��\��)�5$鋂s�~�e���j�}��c�A}4DB�U�hA�^�C��Ć��H��g�W�`	�F"�ِ����� $W�s>�Ļ�K�l3��QN�[t��$��=�c'Z�ɪ���:�5в�e���O��z2���ss��&,����Xh�Y5�e��K�û�������x��<"����� �Ok���f���%�)�:�������v\�x�|]��"~y��Wdi�ھ�騍�x!RH2��U�%��`P:]�L���1�~�ƻܢt���U��u�Z�qfx�����X��h���z��$y� ��kI
��������m25B��
^���I�:<�%��8�c���GI�$�f��I>������H�ĥ�VFCn�`�{w��bu"�eP�Ѩ�1�[���h�X!�~}��s��r.�K=�P�܋���S1���4:�����l����x_�x����J�^�%���r���:�i�e��ú�Ӄ�R롪�t����mx�J/�¼�
�6�����-3zx>����?��,���2s���Y��8<˹�L+�/4
��ɇ�~3V�vw��>Q��:���,J����rg��O_.l�S�X�6�4H(M�Ȳ/��;�4�D�+�觿k��uT�­��	C�;U�A/�T׏�Ҭ�Y	50K'1	����ѕ�+7�B��TN��V)��;�.v#��g��""�+X�MTf=�[��~�Һ�l�x�����k{���'�mU������I�h��<��-tz��$��⎛��=�>@�;���C�����Q�-i4���Hv������fp=������O�ם�%�q�S8�&�_BT.I��/`n��F�Ee��r��wT
$k()�.a�O�R�fU�� �s�j�]��uöj+5�:'�Dx�����D���F/�yQs�zx��x^�J_N�g;��k���[���co|'�A����yW2@&�z� �Y�,$��xBrB>8z�2�䰆�"̠Lk���|��_����ݨA�'vZWM;���PrMEۤWʳ�ٵ�Q��L�<��QAڠ�k��^@$��>��������!C����-��̆?�KQj"#���M���X���2�"�Z@m�Ծ�z�>��C�#�F�L�&2Z���icZ(���a��Z+^K�PR�֑�kK�a�%�#b���~�a���s�$7�P��׻�<��*��q���Y Qr7c�C��g:����kL�A�(? ��m�\�����&e������;L}M��>���II+:(��	������x�<0�h�łmL����̙���8�5�C�ֳb8��:�:��p�M��r������m�a9�v�,���ZcHpU]��I���<�,��M���K�{��M���DGb���(�Eb{=o`��f�#�^�g��	݆�Y�1p��E���E(�{��$]��7�>.��B�c�����`���@�4��i��il~oX-�/S�I�.t)(P�Q�j�T2uy�{9#j�"��`.���/��Y}z�;3����
D��󱬪~����%6e\(�ϭ�l�-)�`\�Y��M������Q��0��>�9��Ui'�3y�$9%/X	����Y��!�1�1������m��OHq3NG8��p�P	u��T�qĉ��`���B!��|T�K0_��˽v>��X������}��OD�g�H�D�6]"A-��h�/Heכݑ�8(6𨌃�J�ό}8���
	$�A���s����n�%�1B�/�3^A�Mc�9�ǉ���M�ި �$omr��-]cׂS�7L@�41��~6D�QƹM&k
xq�����
s�A�(�����q�h�"^D��0���V�9�3�j���XV���mMK���?ml�]����%����=p�[�@1g�S�cq�1�_���Գ�2X�mP
UU8-%ܧ��B�
��#��}w1��Я�`|�����Nu��"[�d��a���o>�
Q��۔��yv�Mԁ� ���(j���	��A~E�ux��IRZ�$��྄�j���ңꬸ⿞vy�h-ٽ��'��wRO'^�#�z$=r�д�	���g>&f�7�y���r���*`�UDCuu�7�����@weG��?�֟c:}/!�s0�[�%��)��.,y�)�-��|.����bY�4�;o�K�2-�,2
�}i�=��*_OV*�n�H�Nc��t�V�F?�/���(����[I��$���F������b�#^�h颌5.����m�j�$x)���'i���f.�ɧbR
P�%ѪPD��#:B�Ŵ�/�Ȟt�3��;0Ex�V1�^���8 ֫�v����{�����?!����l�e4��~v�����Pu�2���mw6�����6����T#p{>cZ8D��w��,oer��Ԛ��m��6��	8��M��鲱�,r	�!Z�Q0=v��#$�m5Ì��,��VK��/f�F��O�{�0ޛT3�$Uɽf��'����9�R^�F�m��Q-��lf�4?^p�%�á;{��jG"�6;zMR�H��L�m��H;[�a����ߠ�MALА�) �6�s���͠�ȖD�������A��έUr�֖^>h-��;�PGImn(����?_G�Y)�Ջ��u�A�%wL�ET`��J�2�=08��W�bf����3���<�W{�`oɲ��R36~��"3B�k����(Z�;��]�kd��G�C�k&���]��M�mF��V�6��e�����P��m�.��t�|FԆ0^��F]z}$���
�|0���U��ax����~���2rH�.jN頤V��}">��y]��#_�yA(@��]��P��id��*!^u��G��q�k;�t_�P�
<��9���|��'�C�r�{��b�|8pB�"o2=� *��^�KF27��R1^z t2XQ�]Y���mQ�
��������@6Ppk���|��1S�E%c�0^F�op�;���}X}��nQ �|�@fL{�کX�m���������}�$�_i�rO�ң�Nt��;e�FX㡢pC(&��Cc�2<!��ؖ�L�Z (�L�ׯ�V�2k�Z��K�ơ�֝>�v}��>�su$,�ԏ��9��+�m��&���a���6���V$�{C���7��^���Nׅ�fD��-��.�
�� �G�:����%���ȴ�0,����M_~���T��KWf�� X�BB[�C�J�g�ئ�#��D���*��u5����|��y���h}�.0��}0���Zѝ����(:�/K&�V�]���h�q�"+��l꙯���.����ƻL�[z9��]�`Bdُ��cx��s!rP���Gc���݂Ӎ��,w�s�¥H0-�78̓�4D�UP��`�xS��6>���.��;��f�R�N)��{־����Iq��'��FT�Q����w�XRK6Qy�]���y�c��10F���>�%�d38�`�$�B0�0�����#ٱ��	}b��#�s*��
أ"_5��Vې4�-�ٵy�b�#�A��b��I��J�u'�A�M0R�@��P�4���T�*=�"RK9��\Β�P�.����]6O�����6$��}�d��=#�DԮ�)�C?ᧃ�@!JV��Ss��_NA�^'�0�h��"�-yGɔf�������+�����]��\X�,�1��V�$�p�g�����3N^H��Zf�� 66;?�,_/M�~�C�D0����`�=ʲ(a��� �(��̚t����y��n�bt�?�T"��V|���>����P��L��z�_�}�Ѩ*�hx��޾�x�3�e����*Py�gd��=P���TI�������z��K@��~�u`��ʁ�
j���kK����fOe��@��z6ˤ�ڐL�}�b����*��e�T9�2�~����PV�'o��[d�U�qpk�⁁-�� �4m���*i����|�y�!�>�T������
e9Z�|�y;�� �7頱k�,T��[.eoŌ�d�L3j9T�(cF��ɞ���ByyC�3����,u`?��ɧ�:�MZ���<���:��SW;�+_�Q�@C?�,lԔ����I4~�=5��2��]�`Zd�N�%���!���^�~h6�.��j�mo�C@

�۾���+,䆵���g��d(��Zh�d����)�xK$��}���K�R����X5$�3>��Ri�8llg��4v{�Rn�R_+G/Pu�#.�t��<ER�1�b���i^3!��תXƗg7(��	/��D(
����E��S-���lu��sZ�-3�@�JS�>xx�k�����@B�hfHۭ�W eRa2�N� ���������A���-�K�"o+H�w����YIƕeDn�Uv�}����0��-Y`ы7��\����[f=�, �v��=�w�~�t�&��P��M*F=n�*�5 ���	<|S�}�)�[᪑Z����V��MOxA- ��� 5�)4O4�R�z��r�U
�+W�;�tv������˝p���l��0v��FCT�>�p��lPLw&�;��g�ܱ|��7̢T������� <sK;_�B���"&[ixH+��d&���wt�c_�k������QԦ���2�ф�o0K���iU([1��[��P>��������D�PJ06��bi�/V�B�Oක_�����z��f6�<!�����I���YW65/�a��T1�R^xϭ�v�Ep"p��ȴr��f��H�{�0�6�6Z=0:>~��.����6��~���ȅj�)T�s*zyM���	#�>�a��4�/��)��,�)Cխ��',�Y��N����I�?Ic����M���A.p���X@��wK�;h�SQZr�P�b�`)I�	H�I[~ۈ��ݴ�݃�O^����t��U����&�i4�ֵ��@����S/��:~����pb[�
*O��>HlN!U.�fFb�o��3�q��5m0�8�S�Ȼ+�2᯻ ���j��G0��onU�����3D"�����`�<���$P����*���]�:��C6	����Ґ�n�l�f���`��|���1��85AI v7�k�574�f���s�R߲��ܷ���R�2��Q��\L�d>�O�~|��Y�yO�X(\�`�NpAe�����*�O���=	9'�)�U|�_rv����\d�;�A��ӚL�7+^�y@]�5�^p�rѾ˱����-S>D��'4s�6�?,����Ө?�[_�^JO����y��p�����Xi�{2����H<bLL�;鈦��D�؍�F᎕�m���t�Ӈ�߄�؎��I򏀯6q抇�0�Dg&-�<��+���t�릤��<4�*Ge��o�IH�k+�jE B6�����#�d9��:�����S �}iQ�E����������^�	�N�.ͯl\�h?(,�^i�*(�w׳��� ��-�&�C�|G&%��l�c�ߪ���o���cڹ����߾pg0-:1���Շ��>؋���f߽+�Y��n�����<-'�잢�B��Cٳ�ehoW.�R���v��@�$� �/�M`�g����҂
���i@q�1� �->p�%�67l�k�$`ך�E�}	�=iZ+�	���7sKn��Pn�!���@%�k��fQ@Z�Z�BG�3�7wzb�9�/����{b��.Cџm�*gW�.u�Ð ����tH�JsxVf��>�T-��ĩxqt"��4��]�ǩ<#]�~MW�zJ��f&�X�`�|ܫ�p�>ɧ�Gϲ���ө��q̋�ȡ����7c�(]��1��F�:�2[�
�ʘ�y���5[�50_z�Þ����ґ
�!(w��=��`�7��OА�7�s�Qa�O��e$!Ǯ5B�*o�t�1��i�/���z�x{G�&�$�+a��LR�\[BwS�L���k�k�P�GG���/��\@�	خ�STP <di�I�xi�W�y.����H�Ћw(�R�B�j7�@"��Tw��b+ΎN��-��
~�Ԇ#��qg+��R)�j�FX���|��oN~[]m��e��Zg{�TZ�%D0(���Aw�{_i؍x�r*o-|$��.�#Z��M4=0����L��fU�TACm+�h��a���|��, ��E-j����4gG1�.�Bj$�bo�dua�;nJYYg$m�WVv���u7��R3�f@_�L'V�e�7�cY��� �������� �fv�z�|j�ݶ�]�D�3��hby7V8
�
1=��¼�lC�����Sr7�����`��0�f��J��tӺy%� _AM�ܻCLv�'���~�iE��7����3�q�h���*�xҘ2�5r�݄�cV>g��6�N4ި�kø��N�'�{Z����,p���*��D������� ���zQ�&3���3�d�l��|K���4����А�Ɋ��=��������Jx�A�R���E=�S��1���EWC��.���Ůߺ���I4_��Om;��P#�kQ@.�~�$�]��=�)ُ���7Gk(Gl�*vqn���B��h෕6�	w̕n(m;��xu0%cp�7$Ldn.2(�C���ETw�|���*��nK����`���M�|��WCb��k��9�K��C�P���a�_;�	�gj�ឣ\�ѹ�tV�>��"e�ԑK��� �m�_)�Yn��̓��_D�Wﶧ���ޮ,}˳Z_�%1BpC��H�C����;���l�u �`�[1�Veu&좐xߩ��J&59�H�s��s��ee�Ti��ΤpH����+E�g�q.T��3윉�y�� �q���_6{He����k#8"u6�qj�lX��I��?�~�(i��T�U���!a���#��Ml-F,�h��^�� ����y�X�T2��^��W�C��9r�f�ˣ� Zi?��/��g}�jjʮ�H��H=�\�U���C-f��P#��K�4���'t)20�5f/�`��y`�V�钞�����(QmV��,sl�1nI�6�
6�) ���O(�ʆ?�C�T���2��Z�������4��C/�d�R��}���U2�Qq�x#����A�
��cBh17��|�-)�^��).x^"�Jcg�¡ϋ2DƁa8.�T�ȅc]��Jf�N�6�zz�P�T�"��x���k�ˆ������˿�V��y?:�~�Fn�&|�xa\Q�>�h(�"r�ѥ��$9�+�'��wԳU��^k�;ǹ����������ש��`�Fv^w�PI~&i>i�A��NԹ9�fJѐG��a�Z\U�*�&���֜�Ά�Z�u/<zcW�V���1�������� ��f�u�J��69ly+f�b1:v�]�=X~�K���:R�f���Zi��=��>��3�^-<͹:�C��O����nV��L8����0.�ȡ��8�/N��+�&�ߦzgH����?m!+ÓW'�:�J�}n O%.K�Q޹͙�Mأ�n�5��|��n˵�.�[�t�� ��9�.�F��}�*Ř&:��%N��3��.�a�آ���<���Ґ$t�PJw�NXF#����P�Ǎh�#��^m�f���?f��ð��O`��ބ]��H�0�NX��T�̀���X��Jh6�b�_CH.�����砐�x��Ǌ]��'���)��M��z����]=�e$s�h�y�D�Y�r6�"���M;4YHl�U�V\�6-���<S��W���-C4����.�8=��9t}j���ŕ71pБ���
$�ө��u��<t�c88tJ R���@~L����K+�tGoAk�F.5���pbB�ݠ��Z��Z8ր+-$�J�0Z0?�g�p�\�W�n7~�?�t��B�R�0��A~]����ܯi�0�(�LƀU�l��VU91i]��_VU��??I�Pq��U�@���SpJ�g��X����A�B�,{��f�V*K5`%k�$��ݷl��"&��W�0*�u������1F�J�s�k�����?$4����Ş�n�O�}/yvߝAs��c+/����R'���6��C	���T�����-�]R�Umĭ]�=2�a@�v!��x-���>=����hT�E�A��c^Dݢa�3�C����t+��V�5���M#:�	ue� c�)m���%Nም��`9&�#�@:�\�U��1z��3f��#1�:���'��/���t�B%�jᙁ⋾�Ԩa�8����8�QL���"s�U�
���)��֞�:$I[Gʀe.�$�ݜ�s�bpA �]�j��@m�#��������ˬ�/^T�%��]t��[�Vb>����h�c�K�+���(��P�������x������Y�[o�|_>;��<oX�$,�&�$����^�i�j��0O6�"�]����&!F��x6�r�(Yq�O�!̂h[e�&$��F�(E�G��abu�ł"��f��$�[�x��N�Ȝ������\�p?�C�U^q�i���I�#}����+�*A��3.s"�AU�P)�Ja&�4Q��� ��M�c�d��Dҙ�E�ɺ�+�{��ľ�:!(�I�t��a�q�O�{u�Į�����x��_1��>�M��n��|�g3�	���O4w�\f	QĲ�T��E^�!��I�m6i���Ϲ�FP��f���9�&�N;��6Jh��H�5��^���'�I}u�](�ڣ+�rI�~�+�
R,��MW��-ro4��Y�e�l	G���ʿ#�X��	��39S��f�,��Qo�-"���_mL5�]�d�z�����w��Ο���1X1��x4y�!�M��mR��d�r�(�5��qr�y�b@�E�%�N-5�eZ���8���k4c�ч�?|q����p!�o��:T�	/�x)�\ �f�y��T��k�9ۢ���|m�]��HP|c�|v��tZM\��e4`X��ˠ�$�a�h!x�;�T��J۹룁��_�N9*_�ۓGʈ��"���?�{����_���Gn+��ε+��HNF�nX�Od�m]2�*im�Q'��[l�ۜ�߿����ީhGB_����|4q�(�O���8X`Z���3�-B�M}��$��D���xQ�?���՟�(�qO�f�!���d���n����"��Նa\멦>���E�"JL4+�dAt�&8!��eD�
��삼����\K�wLNz�q��/{�����8H���֓��H�B�I��Hsz[\vp5KN�N�,W�����b5i^=�W1[��k�m��4�XW��֊A�uy٤�8��P]Ho윀��xK�R�NUݮU�s&�2�T`}.Ie~������|Wo�3�昴��񿅸Կ�e�~�-R�Pj���J���Bu��Qۮ�L�|>��	�co�;�f昩%e�sg9���h��W����n@��v=���2#�wతNl��]4,(��"+��'�����@�aL]1�h/=�nw찞W��T�6ƻ��zF
{�k�a~�Ӵs�)F��;���6�HǼ?a}*�<��]ps`�����FM��JcJ��kV�Ӣkn�β�1M���S��}K>o_SgǷ�r�/�qv�~-G�^����������˸sɕU]�dJ��X����"�Uu�_�ؚd��<Ȗ�����33�D����O�b:ÈC��B��Ӎٔ�қ'Fk��|
D!��xihX��v�,�z?��#�˹~l�����k�� �$�֓�$7�dyL�9��N!�p \������ۘR(�ş��F̊b�.��� ��us�r{�UD�>�-KY�WI-t\8�K�ʔߛB���ɚ�p�J����ڂ/b�����^��}2�=t�[�c��	1�Pt��� Ąr0$����=\ǹ�8с
��I����~���h��T��Kf54����H��ȹT~��)�lFZ���o���u$s/׷]�e@|ݧ+ky����J�)�^�#2�xk�<��a�|�z,��䫈�5��X}.iLo�F��k�?;�L�UU�Y�*�]%/x?�� Kd_`Np��ҍ�@ �E�3�'��.��*��!K�;�e�.��~�x$~O�9��M �>,1�uN�*���!B��$Y�R���k�W}Z���C�ߐ��W��^�E��2_φs���֔�-dI�Q�g���Z+O~������N�e���k��d4�#]�t��d:l����Ʌ���G���������/��&S/��Q%�8BU��+I��~#��um|;�8|�tl�8�|Py��ڶl���gK����,)��V�
7����P8{�#w�ܬSϹ�_�%�a@L�4��1Nc�9�bc�*/�Q�Ҁ�}���F5�Gt��,��B^��}�-�-2}�k�<y�(nO�p 7���O��{�1)58	,�(����6K�	�%d%�������)�@nYdm�A��]��'C�	%��A�D��0�P9tO���ε�2*�W���D9ys[��9�������E�dMi�6�g��cs� >���`"�rM�10�������--_ɻ�(�<&^ǈ��NQa�	�g �'���B�w�"HD�w��HZ�N�U�R���*4-Y>- ��?饒��A0Z��d�⾀�W��՜��'�t�L�B�b�ŕ��x�]ru��C�XJbT}� �Y�O��:"Yj�aK��,�1W8�����}���;��a��Q����-�� g��<
�,�09r��cA��7Q�S�Q�k�g���Gu�?� �����H7����<-pdN��V��S5���L&� 삊�9���W��_�ѷUH� ����_ĕb�ٷ���05x�6P�!�.���4P�6Ɣ����Py!����%��$��M�"��5OE�6�ܖ��@����ߡT�S?%Xj�M�䰋�C��0た5qVMc�$��s��p�w	��<r���?��eؔ/PW�rܓ���Z��Q�)�-���^�+�V��-�d�-�r��w1@�"���i��,������i�i9t��L���	�RER���I����x�9�[�gA[��T�^��8~��8Fxf�9P�+���l��5"C�������F���W���·�C�N���V|�&<�.��^�h�W���1�ϼ�8-�xU�H�w�������c*�ɪ��Go0�ߓ�g�0��`]
�(^ǭUhV�3D���k��̼5�<�2ۑ���V�	@Yv��0���f@k��������Cۤ�������xA����<��c�@��u� �����l�v�9�S޴�8A��N2T���A;-����C��yuf������ӄ�EFD���pĬ���V6d�>�l�?V��R��-�i�2���Tep���T~Y>���l����U�_�4I��R_~�J�
 x��j
�_��:�8�݆�B���Iw��9ƫ<�<��4#U�6����$��,�C[����T>�ߵQl�Xqr[��˒Ĉ�syH�J϶{G#�
�N�|�!�_�K������<���#��j�az��߃P3a �������2�a.�g!j��S��\���]��N�HS:�?�O�W�Ϟ����v��'?4����o�a�D�dH4���&�����+�:�t;Ѷ����Fcf?����L�J�AǴ�Z����t�[�o'�_�����
Y4N�O��D����-�K<�#�y��/(��0�j�`�����M~"�O��X�咋x�N�u� ����B�oN#�-��_Ʋ#�F����W��ƌ�D&�l����b��O�Q���~f��8�x��TF��r� E��v��SP����d݆���<)����o�!�������X�y�햯��.|�?��
�~;[i½#�@߻>Zs,��اwZ�����W�|#����o~"{��U��������I�)U�8>�����A����D�t+��L�+��i����w7ើ簣�8�`�7��
]X嚍F��BŌ��R�A���.�vQ��Ǿ}Y��@$��V7��Կ(�nB(�/�t@`
��Li�:�27`�Wf�:%P��׺��)*���C&�V��J�,�$W��#(ᚎG��=����n��9�}|��\��xNe\"����>!v`a��۶�/�u��I6t�&uiα���"�C:,��|�.��7�W��Or�N\��Nln��i���ɛ��դ]X�/�����ꠊ�kv{f53��ՃP�@*�<6�SJ�`����TO�TuQVB���рS]vw��_�߈DO��A6Վ�p�j��3�%�/pp���=��7�?�d�~�0̜���1[�ج��߶�t�@8-��YW=5'�� �x��Y\�o����Z���@n�)"�c!+��*�h��1����.�Ŋ�זy��O53ǩ��l���g���u\�{A���/P�֏x�B�+�q��7*	��cf�j�?��*��/���\=��Nk�f�|=J��F�����Z-�s��]������E��N�tcn�����$���]���
�\��`��U�ۿհU%Z�Ι��楼+�Xʼza��w����겜[T5��q��rje4^s�&K޷��`�,9�G9��z��r���W��-��	B��u��e�2?E��d].*^����8�����2��nd'mO7������z]��a-*p�P��{�����H����=�q�#X4��HkҼ�a��%����P��go��f�[Wy(#o���?[OI4[6">H���uod�2[{h���\�?>�Ӿ�o.�	��^.�[�y�}������r)io,�s����^\�1�J"^�a4�I����p(�:�=P���.�l&� ��|�X�6�1�����B�����Esռ�YB3��al�G�d�e+��0c��ר�֠M�������0�ցga�y<��}8,��$M�%���+Φ�;�aK�M�sO%�{8��SP,��>�G�S�P��(В����i�l���jc�,�a!�(��HN�Hgc�E'
��oc?�}f ��D֮�+�L9L�rP�yg������¤h�}��*>�8L%7����d{��(
�����{B �>P:�"����>a�aV����������#��ō\q�!����ʞ;whu-�'צ�Y�wq�j��rv �,��G��aG(؅�*��!���Ȋv���C��ћ���B�&ZHO�8&��c���;�;�wЉ	��l}�eڱ_Yc�5����,���⟈V��Z�ՠ��	{�M���C<h�B}L�����$g+8��M�J�;^���
�����^3qq'�:��@!e�"�/?��)�������I�W�l����/��E�6�I����T^�"���qk����r��;��8)iV�9�bTf�V�ϫ��Ze�6d0�/�N;��C�!��o���,����|�kf7�C\&�=���_�u���HQB��P>M��~��ZĬ\���Y|��9vU29��9�N_� c�N�f=�o��aG�(o���#n�^E��|�Ĉ�=��2���	L�ä�G'���)&�Qe��\:^�A��%tpPG��O<p��"\8&�ak(�KG��$�%�e�{�9b�]F�%�~LBwߴ�y[6��eJ��-(L�1�ҍ�Ͻ�Q2��c�}}(PX�}�=t����� H'm�Mm_G��ٞ�&Uds��d.��yJ�[0��ͬ���wO�^�9īv�܇"TH�<2��̫IHJ&~&/K�}���Ĩ�&.��eK�nA)um��Z��=`���$r�N�b���_�ļ�_QQ�~�?�.��jDV!�o�s�:�v�I'���$+���i72\��2_+js����nw��U�����-�!/�(�csL�t��MN0\#�Gt*�x
2�@�|oh��C @&�ZMuv��e`�T�@�.	[� 5�K�$���H��r�E�[Ms�xĕ������W%�^�2���g�y�oT6�����6�����Y�w�g��b���z5��jYi��l�/[U���%gY��}3Y5��y��n� ���+��vL�[�L-4
��Mm��Y��*�	q��y��N�������ɞ?�W������iS�>���{F�n����x)��;�����[��#��g�N���-d*��Zf�P�OYg8b�NT=��<Y�aʻ�A�P�/�-��@�)S'���z܅A���PDs��U&����}�����qZΟ��6��	j��|�9�
E7h��94��r8�M�[�a�#��Qݱ���{�C�oĂeÎ�♾�mWԒ����]�� �V�ſ����1VR.�D�A�ٯMb�Da�%f0���l��4��^�� �j���S�O�F��N����f������v��N�{,^�&���a9b��NW���q@g����5�zЮD�0�i�<�1$�7�}�F-�.�Rm����s��j��'�SI"n5s��,���(�������(����{�Q��R��^-���#���v7�p3s۹�F���s�։6z�1����ߥ.�a�$���83��9�>$S��ha�ÕXe�uͧKn$?oac� /�-m1����c	�����Y���3y�fVEX�F�]8�Q�臮��Ω�����H��ܳ<Sǡ{{@Z���V3�r����G=�k�u�bV
��a% ���Q˙AtP8�Yq�����ڻaw���-@�l����U`�g���uO�ul?�=tq��pF����^Q�+~����iΣ�٬(G��V� ��L6�/Z��е_���gx��ѧf����}m M�=:E�A;� QQC���1[D��R�=���A��=�/�7ϻbd�OlOo�{����	�<���s�ĳ'����o\Ũ���F�%��j���@�������
�/���`�f�����Q<}D�Q� Q�����n��\l�ܧn���V&0Jt�i�2�g�߽�5g�*��b�צ~��=ϗ#ܣ��������q�(�z>�p�OL	��ڭ���ƪ�q����lK9�X��U����>�k�pG�u٤=��� ӄߤ�jq��-zG�j^c�b'4D�m	r���ù�ŷ5M�W��{>�N��PRӲ�3
��O(鼂�VM�rȶ�=��?��cy:�����D"��J� ���l]���7����8A0����>$n,�_�s䋟$�y�g�kG��q��VOgX�
!��R�����iIaa��G��gR��k��[�7Ěy�����47���Yٻ�)�}}�Ԃ؜l(�z�FJ�Mg%�x�Yf��@t��"�}
G���XK�>�l=��-�,��%�W�*���;P^�������\7�G�<@;�@���X{Rг�`�r.�p��ŕ��r�R�ݴ6��l��4���
ץ�z�X�1��L1\�SWG�����U$cT���������dզҸS~��D��^��Jhí�mǤ2=�tU���y��Ŝ,�XNv؝��x�3�xv�&���b�^���aH���+˞p�Y*'odP>,ִ���D� �O���4t��J�\D2˥��#�i���1`޽_M^�hdDcm,�|/��z#Ǯ�X��ԟ���_@eF(�P�i�Shm�{8�n��i)�N�l�a�B����m����@��z��y��d�-6Bg/�pQ������*B�/���Y��چ�B/%m��޸���l���|э�V�B�=\���iį:��m��~
N����|�8eG�E�LK����wNe�4�r�h�B;�%9B$"7ଦ�{"�����dҪ�
3���3)*�������H�#�g�%�ݻ����bE�L�J~k��NDc#�Se��م��������׉69�X�'�״�@�U9�H'`�(��LkL)G����"]eJ7�n�iB̼��P~!b������e��.�}��w6rJ���#�b��O�y�qJ�*Sw�\��S�7�Hj]�}F�!x>V0�_y���������iD?uB���*ں`�y	��~@�yʎ���亱�l �3e魣���ӣT�p��bO3VC?pk=��2O~̝��yص>�	gE'����q�5�7�ǹ�;$GÎ�+;v�!*Y!�i�0�F�Мp9�*�3�F�+k��[�TB�F=���F�Hŋ�?�YqR�����D'0�O�I��Y0z� ���L�1�U-$,ӛA/������oZ}=�F;����k-���$ʖ���YaH�W)��Ų��$��d,�J���T������*�k�F�Lt��D�ۺ� ��U���Q��L��M`���8���B�䩛��%��E?��V��i��+��=9����L�Ģ�g+8ڴ%L�rH ��ƿC
D̯$��*�7;~R�p�}I��_T.ymx� j~������EUE�w�w���3X`6����,|�&:H�ĘG���2���H��n�A���_+�Ȩ��
3�\�"f�ce������#�C���%b�1�.�FpM�?�<g���u@�u������Z�����_oC����7[ ��ٴ�s����O�7���
�("��`�_6��9�b��Qd��C�V�^�4V�orGs9FC.ʬB�WQ$;ң�O�&�\��䇇/���i�0D8o�L�VT&�uZ�q�8������n�W���zt�Io��fj��1��3&|��@�ەţ����o8
$�������q5Ȇ?a��d��:��,AA�3�t�A�Y暂@�
�SRL�F:d3hV��u�0KH���[�#X����u͛f�h�J�SlL]BVf����
������ݺg�у���|l0��������"�p�������׊��C:+sg\6'�锃������+8Hw�3/ˁ��=cz��7�ߓ3x�k��|��-��jV'JZ?�Dً�/p�Ӡ�0��K�vqx$S��[���E��⣥����m�@�%��=�:G�[�rn�D��7=yr�����@�F���R��>5���h�0�s��R��~���b�KQ�]`�f��pu�,��9���U|,��|ݷ{pf��w�.L��6���t��+�����I�����Lp�.����i��9
���pt�U@hɗ[8l�jQք yU����Gx�ڗ��>�R���T.�Af�]J�x�	��s��䬘���&�Z�h8F�k�a�|��/M5�,qW�>{i��z�\����أ�� C,�a��H�L4R?�0���]3Ŭ3��Z&��ѩ��Ĩ0$)`�2{,b�r�t�:^��hz1v�l7iO&���]��UW��v�a�s���>���� ���eJ�뀀��$J��0��RT�$J��x��0�&��!���.���8��'����ϰ����]��^$����DQ3R#���N��[����9Wq�
���fNw�Q��3���㲱i�c@�G�0(���|�f��b�TO���x��X���5���&̆iΰB��P]���5���YN �JkX�'�OPj��C��3+��%V��O㕼�`�s�c\�c���O���@u|�j�/��j��t2�X�@}�ETF��G3것N�ɼ�e7&�+2xL؃Ew�D�:�Ǟ�h�`Sr�Cl�*�l9/)h7���U�_�Z��?�\F�/�{�?�QVvc�P�I���K;�fAw�¯*얽G��H�u�k��IylhD���U"+��?&�$R7�xh�\1����4<&?\���k�!�q��"��.E�Mo�{P�a�,0���K��ݦIGIV��1r-&�.
����;��)KW=ҏ�{^�+��%V�]�L#��Q�>(������K%/�
����$.㥣F�k+����7���Xf�2����6RwqL�9#���P��&��*3�x(�]��Tᵽ��"�]�~��U�IzDނ��vI��4���Su�_lUM�Vŝ�Lǯ��Lnݒ��b��D�U��i[�^m��b�đ��f��M����G�h)�Q�E-��D�E4�Q1 �*����d�xR	ْ�x�H�� D-8��c
mR�0��6ͻL�4�Mq .#My!��&?w0DC�f�~U��Ŀ��w�u�O��#9�S5��ͣm()�s���:�J��/7�񘉍l)pk��(v��Va7n����H�҅I� ,�8F.�����K���\�s�[qz_4�xP��#3Xƺ��H�ޮ�a���}yG�y����	�����wۭ*,���R[X���>�bF*(@�����j�z��/;t��2 �:*�R�ǩ�t>���[&Q�H�[O^�������+\Ҽp�?��0�Gy��VK����,�����%�`��Lz�DbڀF�C��>���%�z#<�+�<�+=��g5wʻ\� [�]���w�K)K9��(��R�������k�Qm����択�V�łܞ1	l�mB���G��U���+af�DS|�Al4�Hl����'�)��ٲa����`W���Aw~�ك�������� c_����,`�&���!T|ƾ�ս����"�Ƚ����7�k��0��No^a�z��HC=�0�h/��)��t�l���LO'�P 2�8���2u����/6C3�/"�FF�,D���S��عn!���7N�8C��a�����9k��}�F\���ը��X
���k��)�2`�`2�o찝I�F�5����	�t��H)fԻ�־�$�|�a}@��["�$�e+�v���x����5C�_��԰��hZ�ʸv���zۙ��	��I��p/��;�fy���＋�t;G�87�s	]'yޡ�{-�t!�KE|��_��6�$8��2sI�����k	[���?��ff�R�}{<S�E-�GZ�TVg����%��E\2bq�w]��(��̢�Ẻ(�f�e�[gHu��@�ߕ����M�'N�8`Fy".�,����l�x8z��әtC��������˝}��/�c[O�'�]�Ѣ$�4U=��247��Ū=��5Ĩ��0�3,ﻔ��a��h#t��(^�-�\;��MsOn�ȋg��ڔ�G�db}�����Vf�(#�YO�&�g\ۥw�jh��E`��n�Ǫi�Jn�V��^���(/�6_�'.t�����p����"�O.5���H��m?� Ȩ5���2W�j	q�i����d�:8N���]<���I�s\�cr�g6��|Pi�2����Q��+["#Va �P6�n:\� �T�U�ȋ"������ĄHJ��OV1�q�⍠C>��NM8]~��pV�4	��Q.��]�}/��d����z��l5���
�Ru0��g��J�[�7�+*p�w�uhҲ�u�S�Y��KG�ho��HW�/��:�h����k}r�}�=�i���%��,�e]E?EDP0o.���t���<�KO�I�T+eU닽�����?`�i�(�sx�+�&q�-~�M
��:X�OS"���6Ak����uf�+{�� ��_�9E�?��.�22Y�l����R<NYRJ2@B��J���s��y��U
�
'E�0r��v�1���J��T���g;L�K�?�%��EOP���v���Gm�����=q^H�A�/ԭe�9�-�:a���;XNg_��� �ә��Pte{������H�
�j�&($��:���e��_�NF���~h
��N�����j
��d�X�<3��vH��7�7����ը^;����X����ӂX�����5_�������V�m|3����#��.G�.a������U�V A��!"e:x�ߔ�H��i��8*+wāZP&�5��˄4:(~%{�h*R��!T�j�̐c~tN��Gʽ��>�����?p�2�+t�.��9>�yX�o1[��z���Ҽ� @VR��2:)cPNӇNwl#U�+p_��֚�2���Wg฿r�ŵk/ ҏ� �SP��Nc+ C�N(�x�.����,pcA���a��t�þ��~�R�1��ʖ���.c�F�����'sV]����%����ύZ�# u��)j}�f"nf���k����\����Ò�(���*2��B�P�o9�mvJ"�NA�#;W~�@�j2�E&��c����F�k"���MCz��r�ؤW�4Y�W�glWh:_[wfz(,�aFv�$}cGL��N��ߌ����s�=G����Y�~�q�8)u��3�\5.���βZ5�c�n��!(��� ѝ��CI�e�<������Mې]"-���Ν���Ti:W;n�J�iv�2���(4�3�AS��~�u�L��lw�|,�8�~�BQ"���m$Tt��C��wM���� C�+���Hm5t:<B�Vt"��#2(ގ��`;�f���K��^n���8'�c���u���j[�:�J?k[�)��R��*s����<C���&�9"�<ص#y��T�������?��N1��x!�K�ߐ�X�J�G�nK�t��&�k�A;��+K��F%�C���m�O��"�B���6���������$�H��i%|����{�a"]���S�V���e$��k�\�-ռ��j��-02|f&Jҙ�n��U�1g�m�[��M���b��l��d����G�=N51*�{�#�8G/����"�'�-xl>),c��R�b���+�D�~|/P�޻�w���VAAT�ٳ�����}`bl�b�̯皛�����x�U�C�Oc�!�K��~�c�й ��������#\�5	4)hY�deBOk����v⿣γK�Q'��;YH���;w��6�	R&d�Wu���)���v�n�R�&_�u:&f��d��w6QG�0�y���	��u)��<N��R*D�BI�����f2~�Z���ۛ�8_���R4u�e�#��8Ki
�b�Q���4[kɇC����ez��#��w��iVp�!��I���4�. ��<��$e�6���r���m������ʅ�s��I�)�K%X�����T+�+�	��P�f�k��i��)�Z����?��nB�kK�WȈz*g _�[�7����.��h���jMY�Yb	34k1�^��9�y�O��e��,��~]]��8C�F�8��?9ݚ��Z��_"`3�;�T����/��e���t� �g�>o?�]��^+�Hn�b۴�u,���\E��̥ۙ�~׽/�H�V��~�-g*��Ӭ4v	���E�N�t==�@kɘQ!w`�he����=)D�g���(�5<A���S�,x?pD��!9��h�?ajd-W=?��eO�7�"�/n�c��na2�rרjH�R�E?�%~GV�D�ѻR�xz2Y>]p�T��䳫�Ǹ�j����"��Ռ�a�G{���y{�t�>�1CZG���E�N��K��F�)]·-%<��-jE�4Ͷh>LBQ��=G��L��5�\��*����������ij:e��o��K�p�(�x斓�<��{�����I��Di˖��r��7.���,F}6��,�Z.���Έ
!{��XH��� �@vE��I�Y�Y�����G�u��k�oMJ��2�*� ��3Pd��薰u�[�ѱ���>)�rUyHi�4�A��^�Բ���ƐRe�U���g_��S.1�K��A16����DPʤ����Q��J���̠����{+���Jl�fX߆5�h97�V���T`�����O%uuZH$\-7¾_��O�S|?����g�H���*�LI��c�x�Y�~�/�?:]��[�I5��p���Ęƒ����.hj��O�r]�@����e�sq�0�Dt �.5�_)#�W�J�26⹬�)$.o�HWd��(�n��	D�=��o��V>�����Л'/�6򃾑)��	3XN��#�����׭ѥq N~��A��,t�8lǀ�!�cTfI�Vů5L�Ow�4E./`DE�϶�Wi��Y׺7���a%F�f�N!��0=��0+J�u�6p�(Txu���d@1[e������
2MK�����^��܅��=%:c�1�ќ����]�s�����5��j��r�b����G��\e��Cےb�����e��d�����(��L�TK Hh�+�G�@M�J�� Β�d�R�����q>��f4����<x���e|�N-n����q'+�'yv��wc����Jxp|��'/�U���1x�6�4GI�%Gan����f�@�vYUy Vvp��̧p������:� ��5\�8��i��Ù���&��,4�w�K���Z��aҴ���s0p�bʗ��.y[���tk]`#��6^1;3�sߎw|�|�ܻ\v��
�^�U��ޱ�[xq��,'5g���c��"V��k�q�����R�)IQ	� 	+�G�l�����:9�OG5�!P�DS0��E���$F��������^�wPz�*�s	��Dm�u��r���)�Q��O�R�/����,9���$p��`u��<`1�:����iqs
������,�v1����h���:I-�=XEv������6!�VgD!�L��k˲Qd�NE�-��讂A:�|WOGx۬�}�������H^�(\���I���8��ۏ��$��XX��Am��oO��@r�q�:��o�P�.��*�_:����^�\|:%u}^��8��7��.	A	��j�����H�����s�ޕhr�#�+ T��7Pxb�X��L�'���"8�J�!���x�H+Z�.~J�����(����;��~�����)o���_���u_We��h���?�SCI��cpn{���$a1��3�}=��=ն	L��>S-��� `�+���@�C��t}d:_O�rƣ�6)�,�z�V��޺f�xZ=H���n���6�dE��?�9o����9�Sw�����d�iW�f8PϮ� �U�{DEE�t?e�oQ�ݵ��(3f�Ɩ*��-g�밋ؼeڶ
�D��=y���tI�l$��u��7x�����m��Wk��q�p��>A.��+E�\S�o�n�U�L�ZqNz��5{��� �&%�Hz 8��c@e����sæ��=LHE���;�'Ӑ�����Kي߿�,]�`�f0�,����_%��9ی�$_[7AL�o%���b�Q��+�4��,N���~���	&X�(=L�P3Y/���Hfi�x�\|��V�[( ȢFy�5�D�BԜ'��#�Sx�X�כ4�K�{�$�s�e�]�gE/^>'xs���r�XZ5�� �&�n�n��a��z	��:�G�8��Cܜ�'I����� m�퓬��I��|b�N�ƃ�O}4�Cº/���sgVyTEBG�Q�'^C�*�M�4��<��(hq���)��#����%6%���"o�h�s�ɱ<#Rl�CIm� �4��d�;`�i��7�e��wg줎(1�v�SKw2�����y'�8��u�)�Q�f�f��f���|#� R�ݕ�_����F/�	%���f�����4����a�_J�d>�ԗ<�1/r��Y�ýCnԦ\.�/��[흞U���
W^�ǵ�vuL������-����c���,1�[������SqI?���Fb�tJ�;��q���@e0�׫`��s��Fd��e��+�\BD5ˀ&�FHp6�u�-e>�W���H�똰�%��Ǵ`�fh�.�(��3U��[,��¿KgPV*Ӥ!�9*H�`�G?�h뀋^G,N�&i���8�1�Z��$��-K�U�y.`	o|SÀLE�]T�_��:d��h����ag���К���k9h��~���O!�~KU�[<0��p���>jq�`�	�f/"91���Dߙix��pؙd!��c��t����dtdi��B�a+=��Wy��V�tWH�q�������:�[YC���9��r��+���/\y%��.˔�Z�"�y�h���o2Y�桒<ߑ;J�Bt�u�Ik�t��id�B�8��"�j삷8����i�y���L�V[���4����ْQ,˸�xL{�[I��p!��jA�o[}y$���퉕$*�d=��.�z�cbz`��(?*b����(��M|�����k��\z�MUV& ��ܷK�ܜf�`O��x�d"��An��DF���1�J)��Gs�BE7���q�d�o��:�����%��n�%�A�벪umK�f����h��b�ek��b�}�CI����>�LF�`�6R��Q�Ù�@��%QW|hD�>��)>5�?�`{k��������_A�y�b�v\Ke�~����!�|���c0��+�^w0�C��>�x�f,�F��~�Tݐ��Lu>B3���:���Cĺe.I�L�H0%U�a���rm��Qx
��������k·�tmޠ�u u�A�d)	�Y�����~R6�Qfr�㽎��hDķ�ȵ6�Eв��Q�D'�ϵ�,Y�{ø��Q��/$�=7Nmƨ�?B'f����)!�e G�uʗ&��W�4L�w��J��@����ne
�?��!��g� ��,k�3�:�~%��eg���űD):J�o���j>����q���F6^�+
'rwj���7��a$1���y[ĥ�g���Ӗ��2�Rd����1L��|`�n��XR����2��FJ�g��D�}c��>�_G��@�P-���x�]g��&��Г�Y�ħ��^��]��}���j��}8��B�M��l�A�Z�Xi�L˫�74p^�@�
�e�=��/Y�Y2o>[�]���Sm�I�Q���l��P��H m���׵��Ϫ�_nm�K�^c���:1��T�ۉ�#�}�����C����}�;�/Y-Px�e��X;�d�<�tď��4k�ԋ�hpY�	XӪ��$��7�6Rƞ,�7�ʡj�Pxٔ&�� �яZ0�I�~EI��*�%U�ӌH^��[:��SI���G��2fF�[M�6�<i3>�X�@z�Cǖ�����N��
0�SJY`Ɩ'��݄4`T]ó�^�"{���áR�0�|?�����*���O5���Gq#u�d�(�P��O�������"4��Pu���tw'�n1���9&{�y9vgҶ=!Ou�A���W��z�X����լ�9FN��G<?#M�\�s��s	k�P�>/Q��(����+:��w�k�l��k�+~�h������Ř*����_\dt�_��|f�d���f~W��%�]*:,�V̹��Ly^m��+�$�y��1S)����.�y�#)z�
w<d_.��;m�br��'B���SH��?Gg��4̫��`�݉�9��h��o�X₪��m -�qFle�~�t�e�>�~1�{�-G@�M�Y5`����&�t���;M�^�i3 �!��ж���n���(�iƽ�ɽ���ML��¬�p�{�ƀ���Lh�_B�F�d;i�2����Ax<5������q�?�H�@Iꃀ�O�.����7�}�	O`��Cϲ�(B���)3���Z̳�@�6C�0i��	2���N�k�ĵ��d@D��?��U$L%S� ��L�7\�@�YJ���$Y_�=ٱnk^�_I��@!&�)�rH]����h�&�-��5����v�k�;�Jq�d5z���[B���P'��B��!eTv.�N.��耽���8Sǖs{�r��uZ0c洄����M&a�HM�ԞG*���u��!A�����to�̵�!�<#�d��>jaڀ�����i^E>�w�)�x��CE�N�k.�c���ex
�<�K���^/��9o��x���N=?TT��ŋ��X���XnTa���`ZH36>�0;G����e����`Ox�vL��J���� 3��L�PpQ|�V�R0�5�Fs��+�}s0����$������B>
��wJd�rdh��*�ﳋ�q����O��w�"�h�~�Y��	���*����hX��yW�h�9���2�`͛@-�����qrJ�s(&�yIr���f�{�S��J��h:�~�X�]ɺݜ�$ٱ�/@�����_ZP��S�R���I��W8�*Zč|����p�j��D�s���Z�M��X�w�q�1X�lֶD��iA� @�Ͱ�
�e������*���.�:�����`2�.B>h6Xl���?A�!��)?���0aմ�;#ZK ��b�8���]c����;����NQ��>1�/8 z��Ft5�E��[�5��f)��\��'x�l�d�$>(��x`��r�����k��;i��x�6?�G���$Ǵx}��d��
W�@�NM�Æ��J�H\��	�tOt-UD�6��a��y�D�5�4��XV����`�^|N����mdϺj��h���/�K'56�@m�Iؓ枹�fY��f6:�aI�I���ī�3�+>�oA�N���2����"A�Wp���h���g�.,fT�9� CG֥6Hϲ.w8��^fd(߰�m�4�ځuJ9��<�X �z6�į���6�- c�z�,�y�)�H_��I��"wg���>�Vi:�Tv��o�
0- u�Ϲ���>=���~Jqh���v;�<)��h6O�k�v�?w�
dI�/��s����m�����^�m2_��H�TO �|�7�V��L!��pY"�P��J@�8م�}���?0T���C����ն%t1	nO)eT ���17]���8�5a%������?X���JlG�����qAcbn�F��ft4V���8�#Z[<ﯸ�ĸ$3,�'xeyO=7�u"�\�Jqm	�q��S�	蹟�,���1�а���m�ybQ6��tEF�W+Px��K��[�H�D��s�
:����v�����a0�"��9j�AZ��Vmә��0���Aޭ�_J�	���u�d�%��������w��R#"1�R���G%0���='���K��)���r���Ϊ)�%�ʰ����~H���8�K��Tg�p�@x2 4"���_}UW��_+��~/�ԋ��W���4�II��xeF�*��uf3��|��c��	��qF@��(��P��՗T�.0/}�q���3�����f�2A���z�h�e,U����]r�o�pnaX b��ԡ8P��A�9Wq4�������H`��o���؟�-�3�!���p��{k�?� j+�Vu�yk
R���xr����u� ?�5�_�_"U���C�I�iX��x�`v��f2��Y���ւnm"ēu�~ �?���K�6) ������ �ęߦO�éX��A��
��8��P�Ok��+����aY)�캮X�G_D�
�>�p���y�@W�[�������z���6�nA>
�������X�ޥ�٣H�R����U�NPl�}}6P$r��Yz��a>/R�kIY�S�Џ�ȋ�����ұ����ą�=�q���Kܣx�����~C��"�Y�r�7�r����6'Şd�n�D�]� ���tC�81��T���Á��6V����_�Q�%������A/��������,$ $��j$�aw�M��7q�b��95��I���Sq��]�Y�iA�����@�HѝJ�%۶Ϣ��0��c����T��aT˕i�I��2������3�J���D�W�W�+[͇1�wY��wiԶ�#�\"��ρ}]Eq����D%�<I������>/^�%� vzns���8�7�]��a�ޟ���fpyĂFa/�+��8n���� ��^9��}��b�AӣYc�b ���u-�V�K�|�v��,⤩}o+}��:R��ZzY�|\l�SK�!J�񻩰nn��V�������A���;d!E_&rPm����=���cT�؛�p+s\�:��H����3��������D�ٶ�	F�OG1T5%�uI�)�3�����[�L��K�p���.�B�n(��Kb`��>H�-Aу>S�����t�Nū#�gG@�2J���3u����Q�����>���v��r���v����3��#�@�e��O7�Y�/v }�_�����\y����U��>���n;�o�dW��釃o�GkDX}dl���6�e/B�%���<h�V9@���˧79B#Ia���t8�Yq�SV 
zb �xNن'�ؿ���󟞠CJ��!��ϐmz60sn���8;���h\��F�;��_,䓡�V��!���w�8��F���I��+6���a�Ig�����#g<-z ��{�T��ug��7�]`tw�ok�_�H BNa�(2\&D���W�Sr-;�G#���X[����]W�+�>�J莣R�د��V��
5W���/��w����^NF�y{�`G��G�4��4B_�LԜ�D�H���w{�s����7���O�#-$zD��cw�J�.u�I��hPw� ����`k�SVHF�<$��5���j��!����$F*B�C��M�[0<�*a��K����vw��i����߇w����۾P�}Y�ثJ�Oើ`^̼�h�[���o�<Ǉ3���_B֚��ק��b�OHHkn�>4�}��|5�D�݌L��xNb�� ��W���G�?ҊXLI�!����1r��D��n�R(*ҝ����p=&9���G�N�8����b��R�ĥ�Y�J��Ǵ	�Rq��iR*ljl}�	�+��-�����!�}(�BZM]4�Ez �,��� ��ܨ02��݀'��Z�p�J���� _���fP�F�!�r�̃�
Æ��|�͔h����hIC���-���q�Q�h�"�\�Qύ�S�F�$R|U��j�-+)�vY�ڦ���7��;��lh�E��6>�������v��+z���~���|�����zW��\`t�G�i��OyA�_���*b� ������{��0�2K�Q�8QL���t<��k�pd��d���T�����5��8� ����2Eq
yD0��TU���Qt
�y\��&��d:�r,�Ԁ$傽�-V;71Z^C�������4���^��ι)���[�#r?)���(,�����6y�!�"��Ivg�0{fr�乺��xXJ:�qgU����E��ł�ZX��A�#�ކz�U�eL��@�����Yv�� EC]�m�Ȕ���F��x4���6v���q����M��3�ZQ�pMt�.�к
H�gO+B6���L���,�e��o @z��Cs�B!��[?�����}]y�m���W���V&���@سD�!D�d�fی6_��@��ȍ����W�6ڐ���H
��)k���y�4�^>���h}�C��$`�ccs��k�S���Q��(��#.ɉ��i+�;�c�#���m���L�A�#!x�-��ꈦ��Oz3��Ο�Q��r����zؤ�Joj�Ep1椹���5�S'<6O����}rE�>����?�}�>�Qf���X�I��P��&�����wM���l������2�L�r9��x[��&��93���Vڗ(Y����2�f<��l�ꋜ������r�*IA�k��w��� ȟ�H���@DB(I��_ ��H�,����E;��Q5��	Em&�ϕ��q$��
)�Ӱge��+� �X������EI��P��:�'B�~(��LX���MZ�n�:��'��Y�c4���Ή�g�K�
䇝�s	#5�?n�6"�:���p�,C
{�]�T$�/58@��YB�Чb|�>r*�v��ULjc����f���_U� �sܗ](�f͓���8���9�������@I_�_6��O8 �t��|b�*��2������8(hv�N�T�E7�ia=p�&\%�62!�%�~ߘv�k:%/���%���Q�����J#���i��-+���x�u�h��!5��{�G�B;�dJ��d�x}�8�ڡ��0y��7Y�z�UN�&m�5���K�:��P�