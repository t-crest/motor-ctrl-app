��/  ���;K�i�~ugF/���^vCa�o�z@Z���_��0pam�������`D����-Phˈf��T�W���c��ߤw�ltD�Z�V�A��~©BFk��C��;0q�q���Ż����t8�8�甀�7M{ҹ�V�.�V+Ԩ(��˲U~�!�]'�� 8��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI���W0�u.M��W|'�p�㤕k?��p����e�������P�u �>)�ѲZ��V����Z�]l䐜�J"3�,�!��2#��)����#�`�^�^���1]{�}�ոDK���˛A�t������߂�[����j�ֵѝ?����vhl�`S�����h�B�"�*c<*M\f$�"D����#�?��H'�>G��2��D��8X��Lm�Bȿ^̩O*�Lfɜc�y47s�Q0!ӌ"���W4���r�g��`=G��(�UY�AZ�!�+0#���b��$�h�l��n[�gg\���$���K��@l����C�*8$�ލ1�4n�U	<tM�W��xƇ"A�d@��[���-����p�3�źh��^����S��C��(��/��fVIz�x�r?�-V\���-��p$t�=�=�ߓm��Y��ܩ�T����fTkՆX��W9�������	
3�Q�NkT����ż�;��V�D,1�PU��(f���t]i.;���oO��W��jK�1l�;���}�b;J� j�ѫ�ʧ��U�9�vd7)�ﱿ'�34W��=�L�8z>cCw�^-O5Q9#���b#|�)}��g#�ȂC,F��|��o��V�7-�^!��R�K9R��.�R:�jHaK����@5-�| ,���IË�C{��EL�9��������ñ~p1���d��8G�2f���