��/  ��� ���$�h���ϟ�c�,=PX����I���t��"CH��w9]��~RB�k�ֵu�$Ԧ��ڻ���K�4S8��V�/H�/�f*q-yr�EZBz�1���2��>�m�m��T��h��|��p&��e�(C������a�7�3����\��9���(2��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�cǖ�x
�Ą��8P:`�((�w���岖�E��
���Y��?!J���j}�i��a�URB�P����ݠ�{%"w6߽����}�(��z�MWs����?�[Ľ�H����Exy�[+WNr�X������<�(;�H"�N�k��X�zN��p�����O��`E!��n�*�h"x�i�p��ZvzS ��>Ms�� ���r�e���v�0W�k먒Ԯm^E��#5�`f�~l7�lS���Ķ�a��bd�)��4{XG�w˚���yCc��*�`=w�Y���9}Ki��挞�WR��P+��ƪ�T�w���a�$0�XB�_G�Z�4'p!�yp9�I�{+�~��Zj۩e�n/���h�,�|vd�	���*;���H����ޚ	u��t��Ɖ�r�H�[�X�{N%1s��b3x� ����J�"�/AI\�_�D��^p���m������������_Z��F�H����$��,S��8HJ����RR�
�S9{�=,A��9h2������Q�(�Dc����%p� �_t��T��BW�?��,Jcn���q]��Ps���b���fx������Z����@x����#�Ď�`��\0�]	EY��Fs��s���Ӹ�$�}S��.�pwΆ@'@X�A;X������#��:w��i�*T3�l���#��#J�m�*+|�Y�>�V����A��K ���[�����uZ,'1&�����"��"�e�� ��&�{o�Gլm��g;�2��h�'e=�jH���)�gh�mny%�󍸐n�I		�WlFgr|�*�e��&V���4��Μ,p�~����"�<�H=A5�P����}s!��36�{���OJ@+7�]��^Ԛ>�P�L�x���*
����h-a�z�g��]��=��M(��b�]�<��k�e-��&��&���I;���Y������_�H���+�׶5�Z���#�ێ�I#�������ǻ�Ӷ5�ح�� Ϙ��Jk�o��?�.<��'��h*��+W�=*܃֓3���*���v�(I���d.��KQ�'��-YK=��8^�������m�ɜ��"Pm�k���$��8nb{���8&J��8�f�\��ura��$����)��C�y������%�V/��^���J�_�x��gNT�������Wk_Y�4�Cm({D\���+���	��>����1�M��]}�l>�X����/CIc�R�p��єf.T����ZW�6�t��Y�@����**ݚ�w��9��v�:	w��Z�� ��`��D�"�H�H	"m	�W�0[�9Җ;��\r1�Jۣ#�!Pu�A�b&�q<F~�J�k�>�k/��-�u�~�'RzH�V.K�)O�N�]����"Qp�����J���wR&���+�Zʚ��k�!??������}J��M����FS���?O3:�]7��s�e�>_e0j�p`��⹃�%��3�౷� �:̏�w�jI<ZV���s�x a�6��LD`I��q�Px5�`lfӄ��@h������Wn�8#� ��:��%
yJ�/�<�ѸO�(�#�Ɯ�ySnv8��x�Ճ���-�o`@���k�"6@��ӭ>�^����.�Fةd~���%�5�=ei��\�T�?q�F?�X���
cҦ�ǋR\��݊/mqq�lL��H'cz�G��ş����?Da$Ds�2KI�P�"�jaj���bQ��.��`9�lv������:�ЃK|	io���6���t3�e�����02��*�b�C��#�Ja��nۏ�5�؁@~u��z����O�l�lͨ�d�O���M���Vg���	�"	�҇< 
�b."�U����rȤ�E^Qd����(7�i�+��S_��=O�>�E�&m��oh�������3��Y_�R�s������Z�Ң�8��%n�H�%�ʰ���#�;�R��ζC$,i�e ���3Nh*|��rt��T��S��-H��r��bĿn���#ϐN���0��(g ќ�&��d@] �ڦ������58���7 0���ߦ��@�#T�`�q �fk��Q|dj]�
�t'ݘ�����Y��.A��K?l���f DZ.lɡ���#���g����3�A��	ҏ��٪u4�A',�r�D��oH�^� �Qˆn�}��x��Z�U��\� [���v�Y� �s t�]��{�<5#�LoT��8�ea�mfq��(����2� �[�t_I�?vը��'�j�^	��ȫ!�)'�\�@��1v�j��3�h[4�d,aa/3$*%LO�Ya;�6=�i��Ǽ,���V[ͣ�����)�N�z����J`�"���*��`��=G)b�y�y�o��ŷkZ�à]Wl2�.�N}���^�������0�-�ڬd���o���-[E����Q�M� r��E�����Om4Q1˖�v�G	��]x����q�{A �L��=���/�
��sʖ6L�|q�YN�k<jz�}�	;yd����L)��gX'��"�%�����3��b�&��͌�Sl��!X
���5��y��Oy��D��	������.�>�eX���/�;i4��ٽ�ӄ=(�dA�QD����{_=.�������Ѷ��K��1ުQ�t��3Q=5�(�+�֪���b6���A��F�H�t7%�m�>���u��v��Z'e^���U ���\�����K�+�Q-��B����m����R�4D�Kڼ-�DB�^=�O�=����Uu�m��gsmP��D�>L�����+^�M8����3�w��1��	�ptwa���Dl��f������>҆���t����P���G�(p{����$|��r�S��݄�8��tOO�*$ԣ����	��y�^PSe@L��[L��ߚݿ>�f��>��G&��#�s�[���-!2���q'�g�T�;ڻ���Ci��8�ǧ��oP�>u�9��k�)8e�����Ms� ����Ǯ*ۓ\"o���(�\,�8�+�?�� ���A�S��e�<�&�3r�rC�>\E
�ܘ�5�DH�%W�h��.���^��P�>u0?cؠ
�
��:E�-�?�[���@x��eoR���y��[��ZBF�{J)�
Htb�(c�hA8h[R�?i/���(���C|>\X�,�px7Ф)!��=Bq�w-�˷�����2���Y$>z�*[&[[���:�Tdj)�B�Z���p8sT�0܄�����|�c�2���?R'�lkKt�8���y+}���p�t�wj��]����v���w��S
�9Q�E��G?���p!�I�b�̞��_���I&A�ɯb3+	�X��ǗO���(3JiG}U��2��vt���Im�sOC�����~�7;���7��eo�Y=n�W�*=c(1�$��~��
�������KŪQ%���2�z����A�qn1wN��9��]�|�_ccߏ@���Hz�Z>ɷr�����$W2�ߊ]1{��uM�䠇�ݳ���rfQQmuM��g� rYfāN�р�)�f���J�<�"���!�~O�8#4��9�nHeq8ٞ������u��ah��(U��I@�/�y˲v�����,�b��z�E��>��+�9f�B�����0G��������n����9}�Y�����[6����ؠʕ|~���� ͌�X������|��U|q��X�"�{En�^0ViA�),����M���k��5�z�>����\D��YU�/��/�"ݎ�Y��'��=פ���p\�i�JXX�\w�bM��[}�?y�%�