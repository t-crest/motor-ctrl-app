��/  ��E騦�Bmrދ�︊Z ����:�"�>�%�G,���z�;��@]?��{Ь������������<%v�6ǧ�
M��!_�v���� �SV��Ʊ�/�����;�Ժ�y�wK�'N�/��ޅՐ���\�ǗCqF���Od� >�l�g��r�|@U�Hf��l,`x�5���=�?�������ٱ�܇b�Ą�(W�h��\@����|ɴ�H]�j���
�#1�S影��Y5d#->tO� %8\�<��B�V,��)����ͯ�����+��zn���;�W7���Ҥ�LnC:����U J`6�V��57ެz�.�ȑ���*��E��~�0p-X�^����n�����erf��5�UV�`��0;>�[��ׯ�A$�Cq����6bD����Cd5\z�h{����̙�@���?�T�˦b%}� : ǜ�A�irS��|���c��c�_�o��.�U���o���+��T$��U�|o��d%`�������z�ҳ�s:}�ɔ�m>I"j�#S��=\}Ì/#��܆�Ʀ�w^):ҸEpzO�C���w���ȑa�π P�u���X��,�u�N���/m"�V�Gl�$5��{�U�Xx��r[���:�Z�)97Y�%����K0�ev�Fc�ν�<'��d���|M$I���SG9���Ż���~y��LVA�i����[9W��n�;�(�ϰv�ɴ��Q�{IWr���N4��.D@��hv�r[2����M��d���+��2�0Ŏ#�V����G���T���N�'�����ĝ�>�ĺج��R��~����V�U�ȶ�8�Z1-z��x�B��1�����	�r(%a�O���� ����w�t�dU0����WfK�4�p6���R3X^�/��񺵅h���s7�(�ݢ�A�%Ńf9b�g�-~ƣ������Q��D��)�vӜ �Q)�|�g�&s�lx�c��:9�~-.�e�w�#�cT�6؝��ߑ��$�S����OP^�Pi#�Wn�Jc���%g�������C]�8�L}�[�a�oTb�޼~,}H�5�Å���W�<���E�]��ڸ=�#�z�֬�Ј
���S4�& ��A������+�nJ/��ѥ�d�L&��^ES57�����9����y�K��8����c>9������@�^�*��g^I���|����g�4)�%bS�5J�0�L��&��Ԩ�D�����{A�/��EB�u�+c�Nh�s�]vN�����}I�x���HÃB��!�7~G��J��sO~H�"4a�LS���=5VOU��H界QC,��j��g"!����yX���1��t�t!>k`x����:-�JU��&[��6d�u�կ��A�}�ʫ��W���N�x�PA��_PMf���Q��o�N���\w�x׻��� ݦf���'��Ȓ|Ȏi�'r�cG��%S��Q��������w��R��r�T��ĕ�K�Q�@	��VǞ|����5����߸��ކ0�}�Tr��|�Z���} ��xa	.BN�����G�����ʨ��w;�
�);�(p�_.�2	,�M4�ƫJ�J�i�Fn�"��v}
� �e_�?E;���U�	�������D^S���ܡ��RW��
�A��
��
�Ke%]G�#�����&�۴��s�O��/:׀�&^����y�Bl
��~�2����/5�ӒE���_�Fξj}U�� ��2�,����x��˶�N�?+?F7�vڠ�7�����^��B{�>I��WS�y�'�f��P��P)OÇ�\'w~
�AZH.���ak�EQ�_˙w���3Z���`��u�B>���}�AC�NB��l�YO���B~YR�c^���X�3�J���W���`l\�1�-��1�ρ�l\�`h����!_��͇9Ey���.8�X�9�v>ԍw'Z��9����Z������������/6c�fw��P�s.;�X���)���]Ft�֭�eR���.�\An� ����mZy�3�"L4�k_�k24y7r�n��9?UV��	O���i^m��J�[0��A�ޮ����m2�
���FŇW�,������4q����F�W�g���ޓ����joT�p�����&����ã>��q*姺X�����%�~��]�sN�8q!3�r�6�9�����j�
�<P�؜}�*l#�j%�C�0�?�����-7�U����1�H�CH�@0��| �E��h>,T�x�vр�p���涛��CK'ұ�s�P�Ī��X���&��,}��u�dU��ܲnvy|t�N�Hi���<�ȇ岦�����?C?����e�TJ��U2Z?\���Bk?i!��de�}{.�!P�� ����5�ĭŀ`#��D֡E�f�g����uU�U�7�m����QjN���t������샏�!h[WV�p4}��dg6ܒ�!�����q�֣N��3�=f��̘8L�*ؒ��%���$#H�q��&�M�*��	-��s�ZT�_|�9r�z� O�x����m��6VD���f��p�U���eX���*�u�X �'�wZ�DX>�Z^�Ea�z1)N���"�9����L��"|���!�|I�i K��Y@�[�YZ��a�y\-w����W@�S[��n�d���}����9c=�~�����%ϯ�S1Ph���&_6{C��1����)��)�����Y� 9��e��0�/�~��9����gbf0�<�g�W����d�����Z�,6K�/w��3�OR�> �m��=�i'J8B����j�wz�]�%H�!n�s^vy�p��J����Ƕ��
ᶼ�+�	�J�[yc=8Z,�Sr�f�c�~�]4΢\#���;1�!��F4	�7����=fmM�x�eB7C�Q����^��30^�рn'��aq�����mrke�ś�� @�:#tv���� ��WҚ�M��N�gY.A���F��A	z��PU�`q7��nۼU6@'�b2�c	pk�a����WEU�ӏOe(�yEs���~��q�.��
"��{7�7�(�:ɢu�sA��q���L΄��5	ܨ~�i'�lٲ6��qvnX�:�Oʇ9�U���Q]̡2o�	Q$�T��.���U+kӹ��Zԏ�~��l	������?J%�:�_�:mt�
�}�a�!�f횘������{�U*��@:ǉ���Q�*$� ��G�6? µmW%��v{�:�{+u~_B(����K|o��)��?�,)��XSLH�>�؉�/�H��<,��\�A����@��c]J�,Ш�s"i�׷�Q��6=�jA�$�����!D�MC:���#�7����霴����d�߶�ns�@b�I���4�r�N�����T��aYW���(�#���i�;~�9M>�eD����!���@l�z�$P8� ����K|z�'�U��g��q�u����H�q� ���<�e�f:���FJ�b��Z����"��X�b���g�[ZL�9��"C$:�b�&cLҊ��r�:�J56����u�⫍�� E/F��2m�<��6a�r�����4$�F��k�J�@�b�\/�N��u�|J�<e����{��!�B���� 9����?I|��Si(g����0��]ڄOR6fu�2 _#�tn+rХ�x��B�i�Ȟ� zN�{ޭ/�C
�H��'lD�8�����0������T���
�9�}���bb�7�ٰ1|�@ћߔL4��O7�A����QԺs:NI�������d�@n���"���;��vz�"�� l�:�(�?��L�E?7+��\;�C��#�;z�g]�tWV1��qq�� 5��q=[ �$��j���rm����n'��k���[�Q���&�ǸG��sv��\��K3�!���$T]�g`
��:`�ST�.��=��(����<)�32��"�a�׵&���{��W�M�:y-��.hMw�-�>ߗa�~@�(��|�V�$X���������n��6���eN��=�Hł#�]�c�w��	[�p=e.*Hc�D�b�Wzr"�a�3i+G��J}Y!�,깮�=-�c�O�p[��3�S���x��x�n�18��e,Q��d�y�uOhm�X���!����EK�M\�O�&�Zb��c���n$˼��51#/ĩ�e��o	��G��b4I��K�d1�wO�0�KO>������U��M����&�	�ӈ{%��9j�&��˻��Q�� %�G��Kao ���j��8G��w�h������ѝ(0��T�qZy�l5�c��� U�b^T6��n��>2�
-�uEM�� n4�|Oy6~z��[�u�)�.��'���`�6�I���,�������JD2�����Ex�m0�~d��h�{(�
���G������i��~2�����U����G�uU`�嘟��:g��MW+��L5��+Нʼ�:������ե��س��ԄEӶ|��Y�+�0�L����<�"�˒4�`<ϖp :�*�'$ϋ�'�蒤o�72�{������#���e�� c|��[!o��UT�UIR��c?D0Ws/K�+��"��������[�5Sb%Ҫw,$^�^��:�f�,�Q߉��%�.2Ȍ�iS�t(�qaL�ᴪFw�Q��@�A�)�.*�H�QS�͹��N|p5��U�/�ƚ%U�a������q8���/@JW3��I�������Y4]&G��N����B�B%t�o.���j­���40�x��e����T�zr�i��:c���ȍZ̈́�,eJܽ� :|����"` +���c<ř7A�>�u�a:���7t���Ȧ8���B&�j�'���Vl���]��#]p^�V�؄j�G��7;�S��f��Dv�T�Ev\��4߆M�QeE$>�Ք��M�Ӂ�anI�Q3�K� =��D ���k�6�(��滫[�X(N�������L�����-�+�PDd~_@�?(��{%�)\����֋�x4Нl���Xۗ.�(��hy���ن�.8���C.q��8 K1llI\�a0�(�������9��=z�)z�N���	�|C9E�E�Gr�S�v��e	y~XMD?�q��0����!�.#0�١c�#����ƜC�8��
1"��'� Bh7��~�.p�3�T%�0��5�5+i8�~D���x�ؓ<�"��:G��AB���Cij��D�5x�`�H�a��#=g�	er��(��B`cݖ�g����j+Q��|�ұ�5IM������܍D>ßb%�g��9&��4����R&������`D��|�\a�VfGɚ��u�m:l�c�t��-��0�/�U�wE~װY?��T`�M�����|����1%Q��`�&k��EN�� z\g��IG��.���2�:)&b��Wz�n,ր�ZU�b�m[KOizL1a9�AtIy�J��D�����
I;M��L�L�g��P80r"-�s6�� �����͎�ŵxЛ֝�Ѿ+z�mU��x���]�~M��.��X5k~qS������+31�y[��<�z�=m�.1n �@�y����oI��Z$��'.�?C����b
��+�%*�����o���?�X�A��r@!}�����;f·kO�Ļ1��\�2g�x�y�3�S0}���.W�-�E�<�������Z3՛�8��c{Y�0��v�;�#��
�a������V��Z�>��%MՅ��M�+�/<�o4�N��j(		zQO�m
��5sz/��L���W Ԁ'kkne���4v\�3h�s瀄�T� ��t\�O	oy�������jÆs�iK�-�Y���4���ީ���;�+.�$��3��G�� K�4�e�z��5\*��7�L&��.tf�-�s�[����� I�LP����|D��p*Ԓ����Y�#k� �v4�1�+̿�k�)޴��ݲ7�W�����y��[�f�x�v�QƑߑU`�����'B�Ck@�jȽD����y��+�3������I��<�jJ���c~�מ+Ӣ���I�ݸ�@�۲o��n�w��������-CVнB#nWsr=�? �����	}���[��A�c�
�� ��y9R ��D�S^�Tѕ�)M�NҚ~P�I�}�1D�ڛ�M+�5�<G1�X��n9��>1[��w�)��~,�T�w�=�_+�I�7���xq���9z�@��(���a���2!�Q�[.�6�+�)�`��IUn�L�>�C��?b��1�fS�t���	�T���RE޳	_�Yw+�G<AWRu&�h�2������r��\ު8�eue�(���\c4c�Fv}���"�ճ�|�iސg�`�	R��̼N������2qAs�,��SV��;ʿ�H������6§�Y��YD��S���6���Hb��&BP����æ�"�~dѕe�u�6F)�^s��,(��'��-�fa�&$��MSv����"��y��r���#v�5��v�I����n�X��V�|����Z�^s�t������3��Ru��#�t"�TM���oi��I�mp��F@&�{���
�՟iu�%��Xm�S?���	?Z�H�R���6z)�/��F�>�M��ץ�4�7���{�!��ט�v��G�7u���4�U]�l�����ϕ���8M���Tk��MA��e��;20���6k͏��$�~�<_��qb2�l��#�Rh3���� (r���ַ���À���YY4	[�	���������~YTcP�	� u�)�Z�\��������%�Ho��^b�z���O,(t�H+���@ �'��#�oj2F��,�x[�t��5�geՈ��j���Q߼lBԁ����X$������J��8�`&�K��p*��{��{���?�E  J�V���%yV2���!� Ӕ��u�T��VB/�s�����i�^?^��YN/7er������=iO��7���ׅ	B�����W�%�~���z�]������q�?���L���£���S���#x=.
˂��J	GwB⹅c"H����i42x˱!��G$���Ҿ�*]���jo�/ǴB�Ҽ�a<"�璌�i��t�RmDC�2���i���Qv~���a�A;Ѝe��!�Fvzp����E&\�X��h�b1�? <�9@�ʔ ����؉�z����	�o�N�������REZ'�*}�Pz��WM���w�$S�XQ彭��.ҢM��ģ/���q���ԣw���NR��AҜ��0;m���)7O)�,<4��gI�^W��_4�ۊa�y��v�Ƿ��}����9�+T��(���Y�
P��w���x��4�[zgy}P=.��z?u��h�vk�ra�#A���A�R+_ l�}���T5׼�	��A����C���u�~��j(�9<#�дp�h���3W�!�\��z�܈S4a�5�#鳩>A�}�ۉ͍�7�=���ZuOg�(!ؠzlw��� 6�|�i ް|�,n�r%H��_V�P/��<�,�Qeb<��,G�V�U5٪n.�-_�Z&,,��|�l�b��=w���3D���b�=oq[�$/u�}���-$�p�X��V�u�%z�DFE��xc�Kxi9*��W�����)���5r֑�|�8�O�|��5^��\q����.7G�f�������_����8`U梅n/���Ի�#��ci����O�G�!Â;R(V$b\7mt�����1d�K 8	�9tc!��rc�܋$>��ߠ���ZЅ,�����Ő:Qk�֙�Y�q�e�C���6�&��rI�i��ҫ+	���#W��j4�h��i��~t)�N��~?獀䱹MNG�&���퇄�@2��¦zR����öb����I�{��ŻO���r=ʇ�Hg\�n�u��CF����l�b�!l����T�<l���,��}=�3VY���0������ql{)�x�G��DmV9)SK�s�(�JP�i�A���������4�1�T�L���A�JMG���L�̀�&'���@M[�`y$梿�Do��4���+$vt�W�\�,2P������p3���"��"ǣ�9쏹�o%�	E���4�L*Gn�`Zs������I�DX �mWEh[L6��B���ˏ����ic_���Vƺݺ7g�e�I�X�ܶ����7h��,�l�@	�/�촣��WF�=w7��BT��Q(K�o�9���?�Qx�\lvV>j .3���ی�O��6���=�E�2��T�]�*1;Wq+�������1��D3�� �S��W�����gHy?������1_�����.�%����C�XkW駥�:́�
��*4w1@s/b	�#�� ���l_%^��]>����řq'��W6�O���ԩ� �1���I���>n=ZJxOjg�L�xұ��&��l�S��a	@y*`���t{�l�ֆR�v�0���mo�m����s�k�2Aj��j�ߙ�:ʑ�a]�ۧ��b/�Z������2N�C_���u�5'����t������oݧ1�'BW&�6&+OUGg�y���a�P٦��~���QDػ��ԋCF2/,�P��xӜo�T�<;]v�������U2z���r޾W{������7�c����n�q�~n�X.8�HL�\v�K[
B��ri<v����)
]�e�F^ ��J�d꼀�Ly�`������yh1�(E���]�RF�)t��!�s��oM��l_�2�`���!et���%4�w�nr�G��}%��j��"*��ǏRb��ki=�<�葆�� QJS�fi�!t<�fы(�L�;V_Pzp����d�x&�Y:���gi�Mu�1оgdu����R�tt�<�n�$v/";�J���"�.|���ɻ?ܴז�7M��%��q�]6M1��@ټ����~��ˊ�q�B�� $}_����#��Dh6�V�&J�=yM���#oڿ�����/	Ԓ�	�_ UX�h��.�8Ÿ���{�w�)�:6�V�fJv	ŕ�T� un`�%�(t�{�cG�%&k�J��t#��}��rǳ��}�̔D� �yx��ʁ��Un�.sv��f�.3K�@qf�̌�7cz�D��X忚�Z�e���rL����L�$	%gv�kn�: #�S�%��)�8H�`�ŴrHP���J� o��# ��m�!�W�Q�1�Zߵ��H�q-I�沅R�؁�oi��r_jõ�^�xZw��_jp@P��ԓ当;˄����r�iuh}�mM	��0o�L�M�)��诘i�~�(�CG��L�I�-F��;O���O0d3�]��a���h�n8BnOg��AjCB?�k��}��4���|�e���V�
ka3�'%6���OΑ�^ ��=�Z���P�
�ݫ�? pj#3Ta�R�,ë?>���񝻙u�1Gw�Z�1�=1�	��\��R	�;�Q/�K�}��w���x:�6�A���PRҘD���[�C���k�&�Р0�0�]��g��%j�1��T��K�D?�i�pF�H����O�jw��n"i�����p��+.<|O��=l-6��y���@+�м;$��a���[1�� ����Y�/(q����8~pϸ�Z,�*�';r�*��e�,6o�R�7���ZI�eK�\�[Z�Ҡ��b����h���5`���~1�(���o>Sǆ�!
���z�7�������׌��"�	���V��æ3�:�(����K �e9��7���B���� 4���������`M�<�Ơ��q��D��iURޖ��9-:�+��)�Ӫ��"gIQ73��"�	�SlN�9��$����A 놖.p�W\%���;O8N|A������D��7��h�a	ά����렬 �Qx;�������	Gl`�"R�2S�B���W�y�[�삕(tˈ�'�$	Ťs��Yx�9�N�v��34F�\����||4�8�1Ǐ1 ��OwƯ�����\r��� H	FM|��I!P٥��ߵdbE�}2Kȥ����N w0��~ax��{0���:�T�\pVW��L��C�i���˺}����9�ñ���i)2��t��v���Һ��1�,���.�K����2&P=���f~_��g�c�I��B�'2�s��f��<!c�o�@������\[�F�	�U��e�x�����9db͟`�o�O�Q��B��3�Y3��S�<����#�9	ou��I} ���c�8�٫M�S�%m�����A��]i�\�tQZ�'��j���4?�'�)��_ρ�~�Cᨓ�%����qDc:�Gx�$d��鹣d�f���d�£�γ�5�z+ّqY�*����F����b�Ӡ��b@�Q�E.p�ғ��|�FYT���jR>���F���S`�� ��w�\o��!��a�>�}�mUZ��`�/r?��ڻa��Ef�C�	4(*p�9EY
c��~`�S=Yz@��DPPdd�F����Gq�Hb}�S���0'�.1��£��ѩ��H��Z��৙,u�B�O&��x�ꞓ�p�н���Vx2uT�'J�\^�*_	��^����`,�A�s��BбfF��; �)���Z��2�ni�]�V-@Xź[p.� ����Ѓ�����m���5�� �q=�R�k�S�
��ꈥ���M$���r�	�շƢ�c�i<{b��n9�D\[M��X[/'�o�ZO! h?��[mp�rP?�%%��{�����}��wlJ(:l��.��
[�u}�:��m�%�c霬w�E�.�8[Ǣ�4U���=�pZ�B1kzm�pS�ʆ��v�*kֵ�%�E��E���(U���:�R�����V�c?�R�1l�F/� :��9-ik��7�B��B"Z�L���β;�Q�p���+7�ܐ��D/NΒ#��G��eM1��{,����E-QZ.�;���|���(�\(0�/�x\|&F*r=X��b�
��&�����& �,�߾�fC&�����Q�Qzk�%II���o��-��}���F���nQ�L�d�U�z����� �`M;��Έ#z�Һ]ۜ��c�j���L�㑺�{�H��-�f�$ʮ�:"Sv�I,�z�|�W/p�����U�F�d�9lѤ�S�ȉ<0[�\���<$ �kU:�H7���ߊ|)ؔHfv�œr�ń���}�P���o�z�`z+�=�����*E29�W��=��qJ�;�껞@F��a�x���J
;l7��=WY����tb_�ʘ�k�׸UJ2�@�r���2�cʞ
����_���w{dEP��R�C���'����Y�L�T�t����32>%� �]�=z���^�������
qL��F���U�Җ�\��b�2��`������Xܴw�� ^��̭9�_�z�#��U��=�J�"������Y���0V�V��-m�UQV�\_\���ɕ8���)7[�/n1��s��@����R�|/\�������d (��FM5�D$�a�ug�����EW*�6�N�[�-H*\$�B�>`�#Wb:��󨔡O��K�ڌh�U�:��\�̢1�R�����<�o,������S�:�R���� ]��u���)mЀ��Q]��[[DJ�~����������������8��Dn����5h���"�5,�L>lu��x�wb<Q؈��������%(a��J�0�,�chEb�hi�c8��]�(���ۀσE�c8We�[nJ/�"���ũaPN�@ņ5�[�n�p���1[�1�;��6 �
Ҩ��F�D��=�L�D˦!j�`\��*�7��묪�{�����G�_�rI�q*O׺�Ӱ��?4��-���*���{��[��8[���l�=P��U0#/�HI��x��c���or@�xx��vdX�6x,MX��N@o�Ý���m;o�),_`�I�Q��0'���-�����iY;7����~n�Dz�>]](���F��jF��[%�78��$��I+$0A�����;A_�sj:D���)(��hc�k�D� �IKi�	#s�����`� #c>S��ٰ8:N���)v���ÈO��1g�_�	(fb�V#D��T�����M5�,�����EH���P�H�����7v�%��`s��)u���T�\%9�f+0	W K��V��	���U�.eo�h��4G_�y���x��ڥx
��M������}�.'��M��+C�o�|�D�уk=n�tO�2N��kI�h�`z���^˖�Ab�mM�v#���e��^�X�D �F]��*7/#�0�+o]�)�S�2u:�4uH���á�$Y�C��;tk�=Ki��x踮���5b�a�8�$�Ղ�e'j0�ر���J��aIbw�ާQ��A+Ju��<��r��K_�ů#S)�KuJ�����njٛLr�X~�PSأu��td�r|�5�� �1�("�&
�㪿P
�Z����{��(섙Op��za�D�a�\�l�2�j�
?���brl6�3&p1���10D}�V�~�3�����c�9�nn�a,8�`�O5W�����qtl�F|˅�`O�-�H�,�g�N��=f�
~h�B�[���|�P\�?��c1�5�.sn�f�!��P�2��k�e���J��7�~��vDF�UF� #��u�����u� ѡd�C>gP����9F`��lO2�i�S��b�J��FS��!�`�(j3��y�0#��|2������%�d����mL�@�b��A|{x#r��ch��������9i�����s9�0�^.u_��=�/g�=���B��kv�ekD����U ��<G�
Y�e@:|�mB����� �ߖ�Ǡ{l�!+�G��mE�ҏ��S1)}���ͦD���f*�E�w۝ٵ�������[d.�QLJA�:�7rM]W]�k��06:�2��,�r�t"�0|?N����<��~���HĹ�rQ!6�j�<�R��� /Kk��5�j±�!�>A���qs���]%���&g�g| �D+�}��T������5|M�D�[�J��RI쇮�h?��e�BaZl�V�ҏ���غ#3�>��af�v�ۿ�{C���歹j͖�	!"؆�tm@w��@�=������m{j�0A@y���h�ہ-����UY,�0|?��|HXБ�ސ�V�ʹu�l�SZ�7(�3��?^#<[�s�.���1RV������"m�B 1�wp�\7!�ó:~p��ф���m��U�z`�w2�Vɐ��P�t���2�����6�T|���j�#��΅r���=J2\���ϫT�!�w���5�d��r���%�WD�A3ӣ�����y�xd;�..[��J���;���h��R�Z�A3��%vIZ���\�)�#�ӧ����tx�In��(�5���
����4U�����`9ԋ�m.�/.2�kp��cNO�˝�#ku�����8o��ؑ����pr]ޜ�$�`g�-�g�Ѝ	_ ķN��S~1��`^����JH���᪹�Z��xR�ŢHA��C�#�4.|gK�zb���2�.ε�c�GS�FG�}�\�y6����y8�<��+ηnG}"�C����.Ҕ�˂��9�Q&6�[�F��7�[./�
��l;M�(wT��]��M�b���X��+ww�{� �W�e�v��f��s��K�]��'M叿�����F��l������¤��uA�S�==�E��y�(�)Z?˯#�՘��A.J��
�0nq��٢7	����X2E�P����K_&�\�\�p�Ͻ X�K��.��l��±)�ID�&D�5����2�
�躂kD�X�z�	�S~ۮ�/E��.z�MA��[o �l�(�?�zD[K�O�2c��&�7?7�~+�/*\M��_E�VH�ݴa�o���D%`�"��'��z���^��8�^��B�������E�ը��8��ә.71�	�	`�_��+Ȗ�� 9�mAG5e�5��'��%&���<�3o{��(�r��Lc��D�X�"�s*K�rօ.��\� ��C�N4qs�1y��Ep�PY�.0�T�"xq�����2��:�I�^�B����Y��*ty���T%���)��Y��Z���6���*��T��90��*��LV�a�sU<�Y��u������%j��e+�W\�_�p^��aƩ<�Uk���6���?�N�!�=���.kԈ�`���V�q(P� Y��B��y�+c'Mq����¥
�)�T�
�.t{*��g>���-�0�J4g��*�q��@�d�q2U�ٵ�c��wo):��Po)��L����Fʯ�OG�s�D��ɅAY�2A��_6��$���G?�C)�\�� ���Y��zoy2N��(x���U�2�w���3�T�B���X�!`��g�oG�)�Q�c���i�
�3�Ao��N��z`G�0�̫~��i�F ��mk>Z�=�l�A�+\Rj� ���������m#\ �7ŦV��n8���8Bs��`1&dx��%</:R.�t*t�8�*s��<2����M�S	��(`�O�Zul?%����.�6�z�8���o��HQ��<X,$��R-[�xfA��+��)a0Jݤ��F��jؤq���e�5@��Tsc���i��?�0��(��S���&�V���7��13P�P�2���8�WlT�E�T�,I{�w��������^�� ���Yv6\ �Up�@�:�tn�ym����x�k>'c7��-$N�6�G�+e?N�a�p^ Ӽ��i� K��M�u|!���Ne?<.��j�B#u�Q����9=�����ܷ�;̪x-�5��a�C���Xz�/0�#B*��?�Z R����q=-YR&{O[쇤6�5�t�y������j�p��"�I4�$+��lXMo�SOO����U���U��F�a�Ơ6<�Fw
da��o*Xn_'�ר�g�M�@^����-�n�*���1�KRv�t��њ�9Y|1����t/Y�/�	ߘ�-���m�A���՗�'~�����:��I���*Y�]���i�n~�z����ŻQWil;<T,�Ѡh�!\�ߧ�d$z�kI��P���H��Z�S�\���@���3�rn'ߔ�8ߑ�܏\�ϗ����KU]�Z^��h>�]�v@]�����<P��x�|�2;4[�ߒŗb|�	X�
�_�tWc�4 ����`���M�o=�6'��a��%�
Tu5�Dz��j#=�7X�\.ё�+�H�ԕ�$h(��vkC�EdL��Đ�G9ן�U��ZR� �Ӵ��G2��|r)�M��jR�K��F��&Y�@�VN�qTm7���j@�Bl�&����j-�L);o/���7S,zTE�~{z*磵?��g0�B���]���0�g�GX���?����=6Lm̭�N�@�X�t�>��;�7�y���a� ���ܪ���@��dV/��?���}�#V^r�(�����X�<sŐV�	�1��K�ŒLl���@���H^��gPXhy�׀Q�n���A�9��9*���	����1����_�D5s̳f�ӝˊ���| @�]Du�d�mԊsw>#�RW��	�|~�ï8�a'MWhm!s���H�"���n���a�v�����{c�n�M��SQ���)2�+ ���W����O5��sr8}S��V�s=�C����]7���8�.���L��AҫQT��u�)t]�I���*q<��s/��uVQy_Z��z��y��ex��S���3�_��<����N�2T���:F<�s������9M�U��W�g�k&Y��@�7"���/��BY��J�m�Q̛�I�E��o,�����	vwx��S��j��|�4z�o8� "(�8sX 7����T��}H,z~�D'v6|I��v�Cޭ�,�h�9Ov}�@`�����k��Q~h�a^%6�,h�Z�Z�<�Ն�KM2����l@��Z	��g_������_t�B��LH����G�b�"d-v�_�f�o�g��^k?y�3���94��~ ��$�PP�ٓSyX�;Hu����ݝ��	�gl@�'+V��n�?M�=wp��G�Z|B-b�ݰ!�u�PQ�]b�fn%�Wd�X�lr!6��_
 �Cx,�v�f��{k�L5"2��>]ç~�D���@0fϊ���u�be ���c�O��@ݳKo^B���k?Cg���
�e}|��>��Lt�2'��ދ<�)�b����3�+RK�w����e����8z�)��P��<�(�g45�Ez�2�A��u��'�L;��:aSp ����&�@z�Q��y��W��q&w���JI2p4�6kV�M�5Ph��-w?����j@R�]�V���X��0���'\��Q�M�#���0z�~v����h�/�6G��`^7��*&�9����£ǰ;5V�c��!��K�ux�=2��ۓt	(WZQ}�:��ԃҗY��<61^�%[�tu;��LlS�[��2>-���x�z�NeI�P�g���|˧��'�|�K��b�B��;|ĭ��� �Ur�׏a��gb���?4��k���Qg��'�a�'c ��,4��w����h۱�;ѭ�O}���{o��V�9Gb`$R�tc7�/��b�W�UC��P�Jr���\}됪��u������q6��TZ�k��<2�
�Q6º��z�j&�3f%�}gUv^ݗ����?�E�o,ܩג;�F�W
������J,N2>*f���YYQ
�U�����;�ܨu^.4�I���� `�K�>9��'Yp���#�`N'��Y^Wy�<����e�:�S#��r�@K���UZ��&4�֒�3X��ش.���ς�ĲK����X&�o^�%^7���49[g\��:��_�|�(�ֹ���g����Κ���#mί�ӽ��T���a+0���q����&<�8�g�>޵�ܠ�G�Y���dG���8��n�MLr�(K�;�ښE����4�f�i@�9���@[|ŏC� H��
|X&��]6f��hE�p 
KT��PL��Yzn1V�g9��B79���*C�I�J�5������K�+�Rnto �F��ߔd7dc�_�%�9r�D�g��k"�9���6O�)L���m-�2��'���g��ik�8����䡔�<?O����2��qhO��Ij�5/�x��4�q}?��I�F��)nXc�P�{�[o���+�մ�^�կ�b<��u��n�	�*֥�Q80۷�`�l@�����_���5��2\�Շ~�2���t������
��B-�X�݀����d0�ͫ�D�a6>��dC��1����@�u1p*]��(Ϟ�D^���9R{�j��!w���#�CE+p�uF��[�^6�CQ��L~�?����3y�,f�D(fb�ѳd��K�t��ڔ�a��WA��T�)3LՄS����2��]O��x�KX^�O�|�E��Ba��e�uA��2E݋3M�T#��<�aA�j��۟��y�bB6�j����c��45I]4X֩K:!��ɷ�H/�e	�.��S�01��I��l�滐�������$�q������p���Ͽ��he5ꗝ�U�!w0��)}�KY�<N� �ak�Dq=����*�ER�9��e�@ַX��H���0��(;��U:P�d�ΛQ .(�e�%4Ϧ��y��b$R�7
 x1�ݭ�b׬v���<��&��w�f*s��y�Ԑ��~����uZ�W�S)�$���tt��e/4e,������b���tG���b/�j!m ECN����M��0�Q�e�������]Ȭ��\v�	�Q�.���Nl�O���<^��ul4�$ V�B�z4���kl ��%�D4�]�"$��~f��+j��'�>���D?_D�ocw�.�2�����T�#��C��j�Y��Դqo4�B�'J���w^�
�g5}�<x
Y�2O`aSb./�	^�:�Q�% �"�m	_���_��4W��yX?x�u
E&�~����v�W��#��,s�@���j��S�6�Ù�m�&���,�ۭ�N�v�/��_ ��K��F�*�2Ǘ�I�&[B�2�I�PJ7Q�J��Qrpl����:#����֤L������5`F�LJ?��?��^� @R��-H�m�E����@5��!�^����K�|9�&��I<��.��&���4��{���;>�C'��Xx(�Nt��Ég���h]��K0�Ɲ ��A���[W����XXz+�Av=���y'�L��1���%����![�b�3e�0AE�Rq
�N	5PU�]��02>�hL�&���IC�_��;
(��#��U�ߩ�EWT�D��I��<:6L�42h7�B���p��nM.b�	H�����偽�`Xt�Sa>e��d��ؘY�`)�@٭k���-�����s揦}�~#�].�J�1
��w&�Զ�l�(�5x��@(Ye�Z��\�>
����ދ]�V�r���&��'l7�m;�v��_����[3$5���2��6�ñ�CW�\OY�^\�%�N�]߹�E|^O�i�]�'�gԟs�j&BV�w)�:� }\��	G>�Hm�N~����Z?�T"%��ƥ�`_�:�a����b�.L���T�g-+Q&���y�XI!���)1�{�(Г�d����,6���!.�A�O��H��F�b7�������u�����FJq8!�wct��;��|�y�"���������-<�>x�!ҏ�x�[�N98�[�|t�!&��4#!O.cK�/R�Gn������� C<�� (,8�{�8h���	�=���/�,����(����<�nzb����S������?^�
S͢�_��
9pћf�4~`P�w��w *�A�𢼏���Deq�ٿ(��'�����Јg���]I �9�I����j����������~W��M���C6���Ԫ��D�ų�i�Q-7c�pi!���l[֛�(y�Wn�ҩee�_
�v�+JRf�F��pt���jG�vS2c�9}繺�Y� 9�MQ�r`rd��>�R��T�/�'�DQ��beq��2�մY;~��کujpIc���)o�����X��$��������B��^��]���ӵ3������J�/H7�k�vw�I6�8B��KQ,	(Y��VFhg_U�"UC������|�B���hB�C�L<Y�)�Y��n���?rF�a��#Aa,�0��n�x�fW���4�~B�ʧ�v%�uME���,� 9�_�#\TH"8��)�Y�,�������=���Ą��`����b�ʔ�^4��4�ޓ���{[�c�iLWN�,�e02RꁡF�|.��O�Jtoay��x��D�Ul����h�R��ށ�(8�WW�U���H�/�ף�N�K¿��-���:��#�G���������v��?R`]p�<�:����'~�#�B}�>ʳ�M:[3r���
��&�E�Z$hEĳ݅���߾(�q gS�B��6�Y|F�P!tO�J�+�ь���(e��r����k�7�	;v:`a6��0܊��U�vB��	d�_���4���H�7mx7��L��@�c�)m�����N����|��|K����y=�v�~�f�S%��@3�V���.���9�����yu����Z�w7Dcr��n)��W� ��j��@��ǣ3u�NRf�,�րZ��*u�,�ֱ��� Lz�;\vi��{��4n���e�H���w�Cג�����l���D-i��O6�(ȑ��`�0& hR�r�����_'��|tѡ��h1a���XTm�<2�*A�~��%؇c���d ����a�$��]j�\<1�2��)�XE�>�bk0Lഌ;(����^6���:�&<@���P�5�
r�� �&�����0��c��鄼�ú՜��.� ^e7���s�K�.Pm�����n�*C��<#n#����{�ț���֌�9,Ww��� /D�3q\�����}}�����a~tI�;և��wޠ8˃��]|��u<��e�j�-����nvS&O�v3� ���|��N��7��Nm�a��RN30�Aύ#7H��������%��V^�O^��zf�|8-�6�-��/����)cv�]L�g�Z؄����j�����XBy���3J|O����!�"j�Y���:�X�5&vL0X��YrFU��^>a��R��˻#>�ZGҟTu�ce�.�r{t��'g��hP(9u��Nx�ڳ
8tEaM�Hz��EW:�^xR�/�d��I���R�
����B5Ȏ�mVs9��#t�����"N#:��=��#k��%�p,��KRɞ&����u�4,�#V���qq�V8m�ܱ����¢�ip��M 	sM����ڋ0�����E�g�6y���X_�2���GL�몹���]��P�h�0�~i�Q�R]gsF��7�����w���7����� r��2�����`tw�NY�s�A,��e��
�� �Z��݂N��ٶy��u��J�,r2�#��oM���m���ؚ	���¤kt�Z�6�? ��l4M�xė��W<1Xp��T��Dz[�?�����*�'OJ�Luh6d��A��!G�t]s)��N���u�(N�yc"�K�Bޠp�C��)b5t^Z��&��<Y�+����p�Q1��s��R���уt`_���4)�1�ptSM�>�xz(��:O���y�+�wf��,eZy�F{5��paŝ��a�� %���	F�_\�/O/��1�F�O��'up̦;�ш�<=�8����yհm���~n!=IM4�T�)�D9�e����}�"M�|��4i�on���f�2��H�x��脼s3Q24H\�`%�f7�\�Y�)��U�j�G2�_����W����z�E�o��R�+��(�Ϲ
����"	b2�$�L�\��8@|�n�1�#&��U3B{�q�؝����G�3>��C�m�'V7��}�m.{�1=�6��@0�(U7�5WI�,���@����z�ke�s�ȉ~mV�$�r�ݤ�S.�IP�ԙ�Y@���b�fdL��R&��	���QO���%�T1����&�Y'�ݼ�U�'��Ξ~wXj��5
�C8Y�a�����iR���j�v�Y[g���-��Lk>_'��9vnU�I;�!p��4�3�O�����j�ʏ�`� rb�c�J�?^���s��h�R}׵��ҳ����_�*4Ag1y�45�k-
�6������i����Zk�q��	�/�O#D����]���iI�]��N>tJ�
�2�4A�vǫ�d��]6:��O"9 �N��MУL�DP�P�6�{�ݗ�rh��w��� b�I +}�9Z��
�7��wB�,�]�E@7�j{1_p�X���<i�B���t�Zϐ�4u�5W�4���j��*}݂Q�j��'�T*�pɾ1��eL6��P8�Gf�C�02�quT_D]�)כ����"�ԟp�b�ٙ��t��N�C�8�̇��hS}dj8�4
\ 19�TCĝ�t��c8J'�ڲD�AMk��O[�QE�a�C7#�DZ;��y[�ys}�u���7�L8����+%SҢՏ9��"	~^ͱ��4j�5�i�,�$C�Cٵ�-hÇ�t�/�ɬ<���>y�Gȁ��������r�pՓ�L���1Sk-l@6ù��B�Wܙy����:]�+�w�����^�e�yN�kQ�4C:
AC	B��^�����d���$ +&c�H匋8�@02�4;8 q{�5��ܣIz��j@P#�\�)'w&zTBDe-�ݟ��{��*��n4J�_��y�f�!�ϖ�+�{�J��w��r�m �R!ִ�p�<��-kud6�������T��j�?������0t�������dg��4��b�"����7�">�Z��5�A��X��ñ���)es�?�����L�_�����T/1��;u���>3AnO1@����:��,3R?��Ue�x~R��!F�	Rk����r��eٚ�ZH���-hZG����^�Z�Į0�#�h:ɷ_�m�=�B&��s1Z�����rn�ս�ɷg�b��t4y+�8�--�fYMR��1@}Y��u��t͓\"ƝT��ieO��O���.��Z�5I@��o��-������$��)�ah���U����I@	���c�P���^Tq��j$���K�ES�����J�+�����V���/�B������+rj|Q�k%)�bY�u?eѥ�8��x�E˺�d�ą�W����#���*1m\x�����U\.�ޞ��Z����Z�3�M�N2Ld����)�aUQ��U�L5�,/�e�A%V����Ӌ��ڇB	��(��Ja�l��X+ѫ���Pt�eĊ�9�0��J�TP�INخn0�n�<-Ln��td_x�s~��)����y)���В�3b!ׯ���
�gcpP��TU��3��14��JsĜ�R�:�0Oa�B�-����:��X�s3�l.�&�O3�O[�Z�Sā��5��s�������54Wɻ�X��Uk�������y���֫U�g)����gXf7$!��	��	B�K�f�Έ	�~jXuA�:	��D���_u�<.�w�|x���hզ|��T肷żRfy�҇TZ)ċ�d�e��z�%�{��ԕ4�Pz�̑�:�Q�}���VlZ�Dv�O��C������=��������p �/����?i��gqxK?�a<������	�e�t�R[��S�K����ϗ�`�3�W���4��hK^����������hۧu*�c�S���J!���u���S���LL�ё�F_��"��0��.R6>|&��o��I4�4'�n���dy�E���J���S�7@���rM:�G׳��cL.���S�[�D��oaRc�>��D'��lK�GGl�\_�%̍��f,�K�~	��(���=z_8o��+�}*��֪��"�B��3O��Hp<��E�J_�xrb�2�:�I�t��Lz�A���|�����O;�h"��D���I]ŝ0�� W���o�ّ20P��V�*�tY�p_^1�!	�ہv�S~�R-�gY��`�g�K��Ly���K��h�"�����<_�B�����}�T�Ѷ�������$/���w�&��1]���)I5S8�WT�BG��up�*r ���MFZ��@l��:wׁs��{�,���Q�6�z%ї���>(�K��.�H���8�w:2_8�v���F�OL�9�̲�
܎��oDi�OLLv�a*���C�q?�F��'��ylv�?��,v�rd�|Hrǅ��)���5/o�ϩ/�6I�c�{)E�cb���L`V���Ј/���&�R��H��ݮx;0�,��%<�Q����ڰ+ЩT�	�u�-�R��#1�A������I���~B�-�X�m�ﾗWʳ�����R�^|��t�jo�<�Xؗ��ح2ȟ� �;����jQѷ�n�Ex�P�5�]�[-�߲8yA��z]#�	Kh�>"G�?��WgB��_`5n��tF]锑'�#�������\���(lv��#wwc�A��`/��$���<�?-����e�A�� ���1�����u|/�8��vC�Ī)�

�P���`��ѫ�q�����U����Yjf:�%�=i�o��L	M��g���+-��d�+'�z?�����G�,WʝO����o��l��%��;�G>���_`��}�P6F`�u�~�֑�H���+>��=� 2���sm:����M/�[<�<R�/�dy��l�e���x��y's�=j鋉�������9��?HI�]an)�����p���
�n-��;�}�oS��v�nH�4
K`x�G�:N3;噂:f�M��\/e���kȌ�(2	�	����i{M
z��9�9�ݒ��>�v�ua*�4�<�����4Q��S��7	ߓR�9W�gY�A��S��� �o3�P��F�*(�XTl��Z�Z��Q?�!k�(��`���8�f�P�I�NLV%�j���Y��ţ{�7<� �B� $^J�&�U���5T4s^W��{��ns�ÿ�Ԥ��!DQ^�T2���d3�ƌJ�.��&?��� 2�*�T�����q��.Yi�f��..J�T^��V��������%��ͦ���)�*�����`4z7�_K�jX�����Φk�6$7X�"��6lD �'�Mꈇ����&&���M�`��!���/}�y;���O��U�*_J�	m��^����bJFv)�Ĵ���>Q ���/�b�y[�1�� Tcv�I@	=YIx*��9ٰB�m�o^0�Z�.FQ�E�F1na����B���	�U.d�V�?U�8�Fm|f���KJ�BĤ�6����|ʬ�f@�۰= J���у��Y� 4�a��X�"����ZNl>t[�-O�nP����y����ͷ!D�v��!Y�Ӭߓ�SD5@�V��B*8�Ku��(�ŘM�(#�w�[nذِt�B1Ix�Nʋ����~50��WR�b��F�G�lX�H��;K������E�?�Na-.d�3�a�����k��@'�}��"_�i�-U1ݗ'����D�G�0��Uo�cUcV��8��?�jq߱�-;&�[�Al�n��q e>�/a黌�6]� ��������A�:�c����aOt"����L������0���8��[	��c�ݪ�m ������w�9p꛹���;E�d�Ԁ��IlhkMV�Io�"8l���y�A��>�{�di��hlb�W�<*I���5��44���V\v���ؽ��m<|.E!�a1�F�inܱ�1ΐ<t.J�N�5!:����E�v0��j�I�Z���m�0�ZT���4[#4��A*A<���^i���<v���%/��|�Y�(�=�a/1�}�`��Е����Q����!�8t�M�x Ve6ED�,;�|���H�8�x+s�牢�Cm`h}p)!��>���ę�/��j��;�?0�e�_:�v��C�B��B�Y�_��`��$e�,b%B�x�m#-�`�m�J*�f����:��cq+G���v>dِ[�2:_Q�n�V�r��n��(��~���xlG�ǘ����$\$�gJ=�%A����Iw���7�M����K.0w�8>��@@'C�Y���A[�YJ���w�*�)3�,	�����y����H�>�x��!ڲ�+[VkL��9�,���.(�"̻>7���&$�o��+��M1�;?-�P��?1�v�S�ڜ���	/�����hڮ�+��q��s�������k�F��v͢\﷦-7q�K�b��e�,}TC�9|͝pd��`C_/Ӑ��Ŋ򆏕��� �`ىV';:Ksơ2��qZ���$ܒ��.�S���'�i�#j�F|��
u���Kw�B����s�Ք|Ц��x�����C����V�-Z.�û�Z8)���ȃXh�Q����-r��ɫ6����1tN��E�g�@c�t���K��>/H�ꕯ���ց�W����rh��uet�XC�z>�8ģ��C�aN�`@�#5`�G���{4�Ekq ��Ӭ ��O8����rң�6!x��<���=��{}7��|7a���0����)�l���s����\��Q��7�����/"I��O��\���*{��[�;t�|B��"�i��N�Hq� ������3����"ߛ�O�MS�@%��*��lDR��ч��^�����S��l�f��2%�$����9<��+����5�Ah��Ċk0�'-'���ecft��|�(������i��ڙACh!�7)�0o%�'dPH2`�) �Ҡ�?���o	g���N��}��#^�7D����CF+�@7����L#\�w�۠foE��n���v�~i�Z����n���E=�m�f�<*3H��G�|A-p�@K��.9��X'Ә}��b9:�ߴh�6�i���:��V-do�J�NJUF#�{��E'5�w6�U˾�>�gQC��ԨtL`�?1 ���v�/2��ᚿ�����y#�~�������M���eFm���Fĭ�.ob�"��*�������`��S3`�3G(F
D�S��o]0���8a�7��Z(�+�N5��;��sj�ʐ�v|X���!��}�����Yh϶e
��E�����>J�ݭ�g�N��U���o��4?�L°��E�BϚ����/(^?{�����s��Zū�v�'����H{�U�l���H����M�F�^��8[��ZP�SR����t�M2Y\��-������i���G��4��8Ĺ���ӄ%_��W�Y6�y&3`����M��B������n��	?u��ۑA#��a�{���[��e�C�s��>��ˍ���-ԅ��g�"[_08�5��ERh��:��D�(�P�R��^ec�A7�Έy�iGj'��$�3j���J�bsFxن:R'7�J&ǣ�����ŀ��o��*�kw	���u�mb��A\+�Q<K�K�>��ݝ1�w�'�� ����~�Q��]�43����<�%mN��<�;��b榚�󸖇�'�����`V��>���N����k��UunD�{gL=�O^�P��t#�	Y]�`dE�A(4�G)�4���^����1��|���T y�1mi,x�Fh��B:0Was@;r�^��~3�^����u�G忀XYI����N ��Jƥ���Ĩ!����xe���ٚ�M{Jv�;�:be2DG"��"�n��]k�I�8�b���R+�vX:sI���^VG�O֖?�Պq�U%�no�b~��)`� -��&�J�%��ţ�d	ꘒ�����~�_�
��k��w�g�.�n� �4t�Nu��q���g�Dmn�XJ�w���]�H���)����`�}5�-�;�U�D�b�ә")���97�����H�9JVo�p��S�����g�O������z}q��%-9!�)���ߌ��_1�r�i��[p�\��qqe_GT��Uc3(l�'�p�w����������T4�ڱ�Gy�x�4`���a�8o/�yZ� �B���9��79Y�}C +��ɽ�6>�o�����i����k�2���B�⮫�z�Q���#���7p��迍v������9Ng�`A�������c�ׄNC�v	%^S�e:)d���'�=��C���f��GBȪ�0�X����C��)�;������Z��M>�H1V�$��f�~�q���w�D��R@���H~�?��=�r��ޜ��>�	zUޚ[Ƞ
Ez ��On�י�W�����YU��^L�!=ϸ�A�A]�T&���>$����z��k���(5.�g��X�q��N;�s|�존��B��0�VT�Nz�����Ǯ��=�����t��Y����E�I���^��)�f,�5�cTs�@2Pt�g_��Kæ�i;
֍�nQ��y��5�?nC~��>ˮ���g�<�K�����ߞ/�����l�x����0��N2�����c�Ѫ���E�5嫽 �	v�/K:)D�b�c7����L�<|�J���~u�q��\��f��!a��������d��u�V�+�-��aiW��.���0V��>�Z�l-�_��	2�$��Gy��	�`��d��N �x���/��z��a9�Ǜ� ۜK
�TNt�KWl14\�f�v$�b��#8Df�����i:8����/�G�G0�#�S�$�1!������/%Mh�7�x���+c�����\��+!�8�1hOz�wV�a�>�㟈l���7FxT�u��􎧙E�&�ew?���"rT��/{�3]�������y�#�����;�~�T�"��q������_��ԑ�/���(������+�1��!
[��[��0�!���U��b\�y�1!��Ӑ
�p�=_8nP:�!��	�H��)%��
^23>�R��u��!�8��D``��\� ����Ȥ�\}��[�?�GZxٽאO
L��0m�%-n�����?�v�����3K����js�>�O�=[OP��;�2":A�>߰��g�j�Χx���EM��[�����~��k*�'P�#���5�D�`�B:B j���pc��ۿ���U·X_��L�nG��߼��g���m+Ӧ�^���/�6��o|��:�3��4�r035�A7Tz]��i�$JI��i_��&�=Ih�i%FdW�2?���	-G�7Ƨ�#wf����WG��^6ۍ��+],^?���O�u	�-��ǥҫ��=)��g�2* ��~),9�&yR�<{��pe�}f��g��\��h�m�r�sT�n#�!��rʑ�T����/mv���M���xԋ��l�(<��0%Tfuf@�=����rm
痫�+T���?��N��g�)������$�(�1S�����5o@�:E�M,t%Sq�Nc���7� 
S+F��6N@:3���e}�qtv���C$6TX��I!r���Xe�(���-x���Y�Ht4�2PFrK�~'U>���_��O4�����T�$
��ss�Ե|� 	�~��oG�4JJ9��,"f���pڪߏأ�	��$q���b����W������2wsw!�;�Z
#�V�4�~ʔ�-#Y/�TD�=�ѳ�zZe�ڹ`f(6j�:��3��[sDZj�����L�J�De'ZˑI-�������ܷ����:	�+�lJ�:��q,�j�!BO��z~�!�D�T�8���XeLy�F@_�󘕖e6iI�Oɼ
��0O���1?zr�������@��|_:_g]��M�R��%�,���i��ag��@_%L%I��_O�C��Q���H�Yĉ�{�7c��O����i�▚�L&=��0l �m��D���,�ʀ��
���~���%���[���"SW\I��P�@��m��<����f�NvI���|�ZeB������?PK��|��.�%��K��\:�qF5bA��c�<��e��\���!�N��I���U���Ό�{�H뷾>+��P�ԬO6�����O��;˿�;���� t��4QY`/���ˊ���P��/��|&J�_3t�r�9�Ie���`�udH�3(H��`;)���it�w�4���;iP}hҾ]�ͣ)���B����Ề�ֽ�>�m(��_R��7)�W��S�������+�o9��$&U�:���Y�yV���ɨb��]�3��&�~�5�U�< �[*;Wr�k����Q���a1n.<5߀WI/�D-�D�mg)�O�/殛��@��%דC�K����˼�][G��IŮN�$������=!F��7
���j�x��k���2VE�����$b�������������z�q��z;��7��8>�-Z������E,dюH\�=��_ɩ�)��J��ə�{�H�h���L���c��
=8{Ă0p�fc���O})�`�{�G�ǳk�O��<P��v��֫��b�
J���E�E4����a	UYʰ�1)5!��m�{�ѫC#�2k
5sC�28�:I�x�E�3����#��VWO|���6=�)�|��;��x�f[�8ˇ��"�{�?�u�]��E�t���l<��|;|�=�j��@^k��(�D�#K���*Z�ā��0�TĤ����9̗YjsQkN�V%n~�x	�	X�xBڲ��2 L�iK��
�q[]���ٕWi�����.��L������6}p$B:�>[jf���
sO&�jNS{�T��OQW��wIя������	�EtH���%{J�n�N굍�T+g
�>����`��*��L���  )_%�e�5�u܏��9�ڄv�׹"Z�dTQ~L,�2[J���Ge�P�
��:c$�0��2�j!������.l�F����|��_#[#;��])J����X�BKM�X�dRu��1P�J�kM�0����w�ʃ��-�ا��r�P~�sG�@����x�m�kG�-DDjD��2陻�������hZ��DgS���Ɩ]`�v��qN���k�	I�F�H���|�:O�*-	v�t�~�%�"zڡiʬ˻�02��O�!�<.0!}���� 6�R�7ٕ�2�d��v�����j�Ű/N��|�����%����1�>n�nc���e�Sf��} �mwB��˕1�g�F@uB��_$��:$��c�iҗ{Ƌ㰧a�Ŧw<C�ʢ.�ڍj�1�K�SI���+8��F$���.�r8ܢ��p��.7��@������{���]!�Ȉ��3��cg���mC����2��j�9�@w�]B�l	�]I;�Te��ْM^ە��7[���|`���65&�l@ (����Ϯ�.n#GV(�L��/īE�mc�cOZ0I}�hr� ��E˛1��x�K�Be�j��t�ڤĞ�c�i�C��XE��iG{q�9@2]��5�.�?�+Q�)X]��CA�{fb�+��m����`Ǫq�&߸w#�1W����H&B���!��\XY�ͅA?d^��^%ÜWY���{�R�?��{���ۥȥ�K䙥:�`���
N��g���AH1Su��1G4C�rzh��E3t��LйBR������8Ӵ5����!�qb��U��/�D"�h��̛,@n|VU �Qt��E�	�>� I匤#�z8:�޽�Y�^���O4�)�}�Zt�+�1qmI`FN�;å�7������`���Ci-������҇��i�,�H��%ڡ�GK)�{�;_��:L?-����=��ޞ��-;ARw��(e6�"+��{���
�ʒ����Y�
=/�<ma_RB����yg��v����+�ټ�ƺD�"a5�݆�xX<�B����i�l��~��_���2�K�񕅼{C�on�¬B��߇wN��?{��7��d��9�Ǚ���pX?l� �G����-m��w�3l�#Jos�YFʂ�Zm엒����<�a<u����A������|15��g%�����Q�L���Au՗,��~L��YW��׊.�C�B�a�·��l�z��T��8C���o�+�󝷆A�kӑ$�S���ݜO�Gq����m�A	44Z���p��Lz���K�t6<�V27��K[��O� ��������>�]�TL�flؖya� ��x]B�sUa���ٮc�ݼ2f�ݡ�)1�P��R�<d��x�M�ڎ�sR�fg��_&eJ���7Kk��&%�̓��O%�]�	x9��O���������V�U����̄��2��hrc���@��e��
���l���о�k(V��_XYop�=ǰ�՘�6�yk�#C��hW,RLdp z�2H���Δ��Tǔ������:po��i���k5��$ټ���X�q����A���P���޲��4�)�a���5���K��z�~1�-B�iO��>҉�f|`��T;�~�>���j��ـ���u(jd�ŋ�\����dbtRPyZX�KQFP������|���\�	�;Sr�A�@NP8%!A@3P��R�������y���_�7�C�b�o+X&��HYS��ׇn�rJ��o����%S�~ �7��m�����3{��-v$~%:��s1��r�Jc�W0���3�&BR9Q��)9��[/��ݐW8���u�|���d�V�6q���t[H8@�_o��X�(x����� ��b���c�1WM�/M�@جؼz)RZ���tm��Gf����)��"
��P㙙 ����)��\��t�j�1�����My�X/R�_����Я�JAd�����_jk�_S�ao�w>�r�0WO�`*l�ᓅ&Iۑ���ua�r�K�e�c��'擉��\�Ү�����x��C��d�O��n_�.�ӹN�ʾ���Kk~-�ά����-��J�8,��GA�\wO�� �kpe���ի�����������Hj����|�&q�q���~���s�ƌ}�S��ÙՕ7��
>d��\��ۥ��"�EZ��B�I��R�K¨z�%���uFl^�H���xݘ5U<Ƥ�k�$~��@h��"�/��z��%�@Ҷ
ISoO��iΒ�Y�DEz;a�Z�N,թd�*h39���\���}���O>��*A��6#��Ed�ʡu�G��u�\���(��W��i~�2�n_S'���ǥ�1��-��ؘԎ�e$���3f�`�
Ѣ�f��a#�����|���c��U������Kꌩ^�&p��zGJ��l'�����ms�x <�>�\G6�WA�z^�P�BY��
�R�I���f`���瀢�m���&�{o#��b�����25Cdh��@�@X��o�95J!���,w��K��0��H8�Ѱ�E�g���)�V�p;�-�vt�:�'�ƈ��Ԍ�l�Y_=�s���CGQhci�1����Bf�U�CG��ڨ��`�[����w�����]���vJ���t@�*�(+?�}��";��ثu;�I�M*���S�:�i��;��P���r��j|i�e��.�?n�t�"x�yÄ�@�$&� ���Yꑋ!`�oNfÂG�cwS��������9�9#�7ä�a��3nrr�xh!�y��t�ك#�~�@�"rUH��c�QF����9yJAz��w
�)P�i6p��͞���a�W��T�������]9w���*�����gb����$^,	/���Ku��|L��Ԟ~�Ǵ�/20�!�k��L�$ht���ԕ��T%�Z������Fl���?��V�Fބ�l�
 �ʥ��h�?e�x���
�ҌA����ho�$�* ��O�:�3�Pur�e�s����Nū�2Y�R�C��V��oN.�cPHay�B,	�6B(��8x�~�T��5�� ���^��V�/�����쉂;�����<� �|�(ꐂB���Xu�Лq���Ďv�4w�c`)%�N�'-3��CQT�7Q�����ļOJ�;��v�Վ��l��n�\L{q�r��]�Wh�I��o�j���a���X���V]؅�
��A����"��SE�Yr/��J�W׾�$Sz��fZ/_����6��Ľ�%|��O
Y�~�f�w��}Q�W�^����	d �����	���×7�P�}�Xڮ���GK�$��k��/�j��nU����ҫ��QJpȷ�	��h�B��xp47�Q�]�A��	��k��ל��Dx�w� ���j��fq���k��^��g^�n��ߨ[�K��^y[&�5��=���u��%6���L'ҊA�k7�T�TM�ľ"�=����CW�\��@`3�ۀK7�RHc�{���e}�V����cYH]!/��Ru;cPEk��\T(o����X��.��gXg&�>�K�0jEOI�+zF�w���.G��q����Ƌ�>ep�"}�48jZ��M�����8w��_��نP��R��@Q.R�z����b��9z��[ �n��b�/*�&N{��'�`7D��8�s��W����׎[ݑܷ4,��ߝr��/V{y6���4bSWx|w��@�qm��^o��U����9�\w�
��}�e�K��4^���/����p!;�öU}�R��H�ʛ	�mZ%I�(�n�y��H��^��t�m�Afl!�O�9���* R� b�f��]��F��C�)�	���r�Ǿ/vyE��Y�{b"k��<�#��0��"�->}�"�����>��6"S�j���Yڋ���ƫ���	XU��6r_5fg;j��+L�z �c_�<��t^�R{λ���"����:�D��	�����.��hQ�eN���+����5��/wc�����SIC%��G��+�=�b��]=x��:c��_��U/kѹ�jxv��Z�?����U�����`ٚ I��'��t�@s9��7u_�ο���N����Q���5�WK&�jE7�0d�}�ض��m�_5x�GG��q�癄l��+yܖQ�E�Z�^~�__ܼe�/�oΜb��;��X��3	��s�����$��.�Y�)����$��ċXp����S�d[�x�󃔜�j&p�R�"�N�p��MI�W	B�
h��e	u�� �S�Ձ6�pG�w�V����q���o؎Y��i�f�TU�sR�{$��N+#,n��.� �R�%����J�>2��ŗ6a6��9'�W����|9��5�,Kq\Ɍ����R��ř��`a����W �G)b
T��-mO�$H4���ܸ9+��$&���
����.Oh5�;����$'&��N�t웠B�߂YM|>��ج�|���dB�$Xr9�v�u�:���x
��K����pu�إ�~</�8�͐�)�-AX}=Ԏ�`�ʹ 6Q)�P aנEs08���=f4�@�VU�7���)��}d�*"��ѩ��'�UR*�?I�
b�dd�8��ٝqL�6;Yz�d������6ʩx}8�K�u7]�ʱ�P$��M>�B4?�U�0�k�Μ���y��WN���H*��wbc�z+⩋�F��ӔzR�l�geb<��l�[�w<]�}��Q�����վ٢/aVu�_���߀�lX\宺<����w�j�v�P҅E�H�ɧ,ZV|x_��\/�Vg�祐�M��x/�R�1�"��e�@%��/$t��� �Z�䈜�o�%<��9l��}q3�q�`�\�h��<k�oH�PX�Bi+�N�h��Xz���>��C�)���YHζMW��{��bw���ܭ%%&ya$�Y|/$���p�'=�0R��$�9h�9��U�d�p�<l��C$�-/�)����t�7y(.��6�<���uq�ڊ����#�4��Q�ZS%C���C�๩bi�a�X�ӟ�Z�E�i��$p�ze�,ܷ�T��ؐ��5`t�g��T1��A��2?\/��ڛ��99{�����7�d͖�f ���x*�`E�Rօ��m�R�b���ԧ,z������ܻ���ʒ�L��?s*=
)}�Ҡ����\%'���^�{���ҕ R��f�S����%P�S�S����1���h���?F`C�5��aj�
�P̉ߏv��:���>�sf�zo!��"�V����0���v4N��Z�r�1�V�]��[��r�~��!;�-�a[n@|Y�t����4H@$ lĠL��h0����*�S~L���"�ŅɈ����!��]��jX�e#���:��Y�b%1�ܭ�5C9[��hE�!��'��'�����{j���X�����s�L���%�g��\��@���/@� �Ij͎���2��Dy��?<xL�\����t2,٠�I��R���_�n��M��|����D>�nKH�l;!��(���FϤq��}o  �
���cW�!eI�U���Ӎ=X�H���n�������T�(�갆��C����" &�k�	Y֡Cr��.Q�7��)�ͫ��7�˚�������[ħ�bcQ�yI�`�pd2x�>=$\G0E�{ ����y��	��"á$��{k�T׶�r���	�g]�3���6�Ihd8-'�A��\y#��N�>�_���\zeq�Dg��C�&�c�fƪp|��z_Ww��\�g�5��A�l/�1Cs.Do#���>׫�@TQ9��h0�z%��W��������H.���:��-�S��+����9XibkCj��
!���C�M��8�,D=�����VpǁTqqj*c`���	���6��	o,�^�qq���o-�4tk�8�mq�1�jU�Ϻ�.��K�Wa���I8��% �8�C�����D�{���jZ4�x����^�X�o4�XH�,���c�x�R?�x�t�Ç�AA���0@7�ĸn���a���v�ۋ7��S�~?h���>�s���]���^��w��l�odx��`���Ȍ����xd��J�c�<l�&�vt���ђֺ����=���h{��TvϢ��7b�"��)/�i{[�z��դ��4.C��Iɵ�f|��т��|:�e�t:�<eUYl�'�"���)��+���p����׌6G� &º��o��]�h���[�\?����T�ֲx�����	RgumΉ�Xy�?�s��Tr��L�' ]M����o,��'�EC��i�Fbd�(�22]���fM�üu>����e��:� N���:YNť��ҟ<�G����2�6H`���z���mQ�KC�W��ų��{������Ո�G�F�YJ����i�n�%�xw@B3���]�oi����K���é��RGi�H���,�H�U6"�<�.H��@������J���:>E��F���?g�k�U	�Jݫ�1&Y�0׽�8|�Q���"%l�1��	򀿳՚Z
���L�߬L��T)�a����]���l�v*�.w��3�-خf#��<e!�*���m�0Yi�H&X=ڂ5y��@���T�y���XB�o`��e��zðY�Ǣ��d��v8��&x�UJ���f��jaH_��eI�K��R����ɼ$4{ȕbt;�r���7��O ��Cld}��;��1O#���=R��6b���a��|���z<��C�k���J��TH�GS��y�[p�$���˻���x"ں�G�֠F�`ӥ�
�Q�.�{�&~D��1���T�
�Ni#���~Z6~��G��ˉ"п�t����4���=�\��	ݛ��X�@9I�x��J�c4�(D�E�FJi8���7��rF��>n�]�VN�/�id`L�Q�I�6�	 ������iƠi��G�^�L$C6�Vc2�S3�����g����`񼣊s�kD�.�NK�n\J��o��qVaN�NM+Wז%f�@A$��Q؃{���6_��2/�,겚r/���T��n�Y� ~�-`5C#<�E��3�)����T��	��̥����l�N?��C ?����ǅ)PI��"����7I'eKJ���ҷ�
��'�[z���s%5"�Ě4mC.������l]��;�m|���y�������.>��׎ k���֟�����&X˂ʘ@�xY0mo�O��Y�8(#=���/�t�rǰ��D�w��n˰���%� b~�v�ӲR��i���,�6xAb�|��Ϡ�.X���{�i�[+�id�xi�\QM�Ƶ�D1���E�'������$L��
�(�9Kq�"ͬwo����!�8&�l� �C��KX�f1�7�,�3i�t�և�A�>������߉� ې~"��m(VD��8.��x��MT�$���W�7����F��
y򋄞` ����y�B�w���!a�yMst�H���иj�<���E���r��>t�M%�~��ꁀ�=V��<VE�,��=:#f�Zuj�4L��qa�:P�	7����o%��+��PO��_��M�
�,S5�%�^o���X�UC�h&��v�GXv��`��ve�M�}Bs--G�7�>��&�ߣ����*B�to��4b�Q*���o�F̍�N/����ۊ)���Ǝ��D��(Vvf���Q?=���Ӆ��6�����6f��L�mO1���)[ ��˻Մ��Ę���2/#*߲�`Z������S4Bw�K{� � k�P�_!�,2����7���l�8�t&�V?�#k8-�d�l�����a�JŰ/�鉷m���� �Mn�~�`�����y5Xh,���4F�(W�!]Cz��0�V��������%NQ���|�e�g0�x��l���}�^�m���0[����K$G�J�r���;y�ȓ��Y��3fϛ���T[3>�Қ��j�y���>�)�f���զ'ʟm ͘ШT�����S^�02\����g�ɺ��C��Rq�~��i��о $j.�0�[��~�áp�KHKPH���szb�Մ_>��~5�W�}m7��*��!D�/W����ʄ�
��4���K����06^�ً|[���.�ӵf+���0��?$�����j�5"m��R���0=9��!z���X��b �}��X�t��L���[��o��l<�t �-
�X"
p����r��h�k�j���ұ�7ֳIЪ�<�ܒ�����:J7�1�Tu/�� _�M��1E�Z��_V��mF��˧Es�B)�������A�Rä˚�8��g:��D ��_T��rd���^��i���]�� w�ҟ^��[� �� XXV��X��� ��'���8q�����5�8��)�ԥ3?���+��w��ɵyP�VnztU����o�G��iy)�2�e*��	�_ @������'*�u�)D$��w��^��	�h%�H��b��%�m1�Z�v~Dum�; �^D>��~�˗*ͽ���&�`9��3>��T�2Nl� +}�*n�49��8��H���>z�޵�m%��<*��8L��Iȭ��%�r�#��d����LJJ�a���"��y3z7C�٦�.�h�=q��Y��Qkz��k��\��s���&M��ْ��11V����z���1?b�g*�����ǎ����0��{^������k��t�#��h��#ɪ��G�	.6n�5?pk��о�U�<'�����5L��4�8��e�"R�p{�+\?ǢR�=ֻ���0�=�v�:��D�lى�Գ��|��%7ZF��A�A�j��k����`* ��wN����������N���X�]b����qأ)�K9���2�E
��p�w���@Ŋd��E.,=��W�6T�|������[fy��7��NVH�$�k�W���DR9l{ �#ma��n�?�5v�!!TlZ)-�7FN�2fڥԻ��,M�c!ֳ!C|5���  7X*�՞q��{�h���CKV-���D�f�%�<�		�Ku����Y&w����yS,�t2���O�j���_����vD���pVV�LUGz��{OW�C��9���6��� QW�D����}:қoI�����7.;������%|���$��\�=�d:v��tI1.����Z1V_e��~�jVK�ܵ�W����_jHi�	�~g������*!�/�$�۵�ӿ�˶L,��P��cY61��l+ �G�E�ޣ�T7]����oqɟ�0�t�����΁��+4��p=���[����/�� �@:��-�ä]�D0ӢL���S��f�n\��jB}���?�+VwFԞ}�\����y�E��1O�+��F��;���BqL&��O��j���5���r�Y�y���5g~{f<�<�ʜ��]Q]�[u@!ƹ�PL��5R�$���+(^!�"�MN����P���ܛ�p�Q����.�Dt!�8x8A/tS��j#(�.���K^��ǰ^��J9�ۣ+̽5i�TZPA�L�	�5Nȶ�Vv����;�*�	��&lN��}�f���i�K��]_�O�O�>]�\��,�-�z���x�Z]�$¯��%�	�<�Gk����>�O�@7|������L�cCR89s8,�ɕ�nw�sB�p%8cu���1H�3 S	��rms��T�.�3x�~��9|�s��m�k��g�ŋuYŔ�M��G��"����R����^A�2��3|w�{��r�/-�"��{Y:՗�,CO�gi뻘��}����\�{1�~ڍ��o\�ړ	 �(�+@�|��x��ZS��h�5�L\A1C�}�G~�p/��ܳ�/��N�[�G�⫥�R[�uG�����$��\DyR��<�L�߉x��� 2���1	q�ȑطϊ-l�wP�"�#�j�NǄ�>A|�2W��^�x��������/��*E$���+�<���Nw1�f�{[�
�\�%����Cb�-	�ˢ%!�������'��aU�L5��2RA`ֵ���z�	�cvbF�<����7N��F��t�ڊӮ�\{�!� �'�i<�ˍ�E���<vY��B���P쎟T�K��1�Ī��Љ�Av �`�z������h�2u��>�\r��4G���I�Y�xX��b���{*�j#ﳐޖ���=�#p;R�]~�7�ʑM<`D{�=����'�u�li�:�����A�4�8M�Z���J�jU4�E��0�E�bn1�K�"��D�� !?�ԤhIL3?z)Ȳ�}+���D��e�|��c�i�}o����@`}�#V8B��ش�ХH��~�Ec�#u�������kZ {d0�W�|o`�s�e��=t�� �Ekۙ�h�6}�tӂe?�Ӊs����F�y�w���"@�&<R�Ǜ{h3��Y��8O��Sʠ,�x���)X�̢�"�T������@[~��>����|����`�vi;)��g�����펴~!�Wa#��T>±�u���_)��wwF
��V��� E������R[p�T�7�O>��䎿��?�a�ێ����JY`��CS	\4���шV8&:Y̙p�.IgT���e`E�tiqj	����'^�-�v�m%a�n��yx��|F�~
Qj?���P=h/�æj�TS�ݢ�5U.g�>��?��55�}{�U�{Q�f�x��lK���eR� ���ﳌ���2J-t�KŁ�'��釣��k`JK��3E���P�k��JwJ��Qp���L���Z �=}�G��3-/��w 3p���W��Q�
���D��$,��V���r���D�	��!{.5��Y߭h�����u�1;/�t	��C$��KDD���"+c(�yF*0N`��zQg�`��H\z �'Q*��,��ko�c8����՝o~��3���S��њ�O�5%qh��[���cx�`~�}����C}�*M7�k&  �g�b����}mܝ\��k���?�^�����u��Kqڦ��lI��+���(t���������M�t����X>��-���,_x���:D͛2|pHu�َ��w��_���3*^�Z��p��3<5�_䋟).���Z������>���~5z����7��������9-����d��CFқm�:,�6:Q	��i+k8�{9��s���d�%���DX�0z�O]����@0���[�Jl��=��>�R ܮ��I/?'��Mi���:Ў/_%GwC��)�D�p渇Ɨ�N|z`��'!�O����Gͣ�n���I��U�����%<L�3`���b�n�v����J��l�}��~N�
����;��?x?���s��H�)J�:0����J�Ǫ^��go��Gϰ��p_p��:��
�7��u^�۩֯�l5���5a��[Ą���3��Z�^�Fj���pN$�L����A�Դ��+�H&�@��\�>H��w�O��*��&�~ؖ2��_����I����JsG�� nګ�8�Ս��,jh}�~O�������s'Q�"
�5���ʕm'��J���i��Y L4��h��y,��`���\�Y+]x� �Fyn$%)�w��j\+۴���i^ٴo�W��#\��3��#PW�5�Pm��O�pȕn�^���-�kͳ�d$�b�t�3�>�r��n�|�y���5�bٽ̖���-��Ί���(�J��&��p�ǡ=L��N�Y9"��^��0۽o;n}L�B���>3���>$SH��r�Rv(�܀�����7����A�"\Bv�>{��J<y��6蹷��i�0e̕������uq�Fc�7;��Ig�Ly��yJ�����u8ČL�|Z;/�jF���-;R�IPR7\Mv�G�/ r�+��gE^x`ǟv SO��n%�{I���4�Z�<o�2kbn >�+^�W]���h�q� � as�u~�60��F���L���j�/ϞV�[����b�Z�A%�-� N�4v�H���U�k�n`��L�ߊ��G���E���9H9���4�߾�gֲ�.~�%�wz߸`r9AG�W���IM���g�fr�9{m�:k��w��>6����y��8�������8X@"�y+&� [XD8��̹aL�\lz�
��w��8�u}����{z�hZ�7��^#�.-����_�ф(U�����W!v�������k���+M*+FRD�¸7p0���;%Î���y�?P�r�� �%MM�O(��^�,��b�tc�G���k;�_$6�ξ46��V�/D�:x+�9qVoNKgu���"�2�(��~w^�F������õ��k���ѓ�bID��N������f�C����ۖ
f�A�Eڈ,��;���4&��',Xȿ	c� �������<8�E-s�0�k/��}��#��˾��r��V���+L������GEh3>�0�i�W�]�k�y?>UKp_�,��9�m�#6*�%��{�ߘ�4��X�|͗���8:V��#��Xg������B��v�z	�KJ6�L�y��6�%X�+�F�^bWwl�'�ҵ�3��CM���b�NTU��y�4|��;�y���i$ap��+��F�,Dx�<�5/:�m�i0��8Ma�ˢ���[t�����5�n�^FFeK�(�hQڭ����x
� ����z;�Ze�cl��:�~;��c�8�s\�:�o��Rx���쌂���V=V{��}|�d�b��/#;~ x$�4'�k< t�� '|��c8	B\P�d\P �{��a�m�T"�4Q��˸�[��Du������x����cor�|����l�i-��������$D�y�^ŝۂ/�)=
\�>�+��4G�x�߫���E�]�{��a݋l�����!quo��6̆i��Γ'0m�_�V�����h�n��W�B�unV�H7uȯ�I�d�6M�a�Lƒ���4� ڇ�xG��9�pXdT���u�a��D��Vy����!<��*X>��z�T�٥�kk�7 [��DR5�0�I%4��p���u�A	�C������B\ZIK1���3O�/����^k�vO�d�3U�[$d˩����[Ƌ�p�e��u��1a��5���
]�[%�]k�;�%]��<ԫ�%�3ǒ���M�HP�~.��֐GE�*�k�>%��y�(�����f���NZ�{G?��A;�߼7!�9��+G[�$bG��돒0�{�O���E����[;h4y�A��B�$"O�"]簑�^�Tm�1�s�dp��bK��: zl��yC<RL�8p2ݫi�8���(x�g�pY I_��̽2����kr��D���>�6/[��D3��^fc�^�oa�ȏ�u+���GZR�Lq֠�E�Cz�z����og�+����2$��&��C<� �Z������X=�D��UY4��Jv�