��/  ���TCq��?��@�Ī傝�j���WD�ZU�D��A�MS��Wˍ�`���.N�݅������Of�|EʅhD��}I�+��'I������*�v�<J�6Z���2�r�� XB��h�PgP�`����P`Âۧ��~{�y��F~��p�+��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<�Rxa?���l��s�px�u�Τje�E2mR�Hl^޿<_���eqی�o��sL<k�?E�u@D�A��(��k��1�	-m:��3�y�8ف�V��]��[=k��VH䅋©@٠yɠ輦V��i�|\%ˣqDf!ӃeӼ�X� �,N*s6H|�����G� 6�Z�`�J���C�:�8���R��s��\���2�.�iAȠ�ҏP��ƣn�b�\��k���y��$ec<��V,�k�ٍ����o�*��u��!�9SΚ�muf����ǅ��`���*y�0�Z I������@���Vx���"i^��>��rqx��,G.�BÅ �V-o��֎_z$׆��)2Ɇ���Z��B�V���4p#�;�ܓ$��4����5)O�ԯ��$�`j^��aV����ߖҝ@��M�*$���T;�ҍ��ͻcu[����͛��Y��_"�?����Z̀�����ht0W�W돠k-
e�������T�f�A�����]�����#h]"!�h�����遺��T�j}���Gq*��
���؋��k��|�*<h��	b�S�1{�bz�?頬��5��kW}�:_�x�m<� E�~���{.�0��7���]
��_w��a��,�,��0yӦ����"%�\�b�d=*ܘ4�Z����k���Pm՜����q�ZM� u:�g��m�ꧬ�����f�W��0F�
��g�-!�w=/���P%��ft���ն߶g���������!�������{��5soBXDsfTx
��x���Đ-V�r~9��H���R.��k�����g��;�و��%0<�.��p^�ĉlψ�b�T�Gn��$�pV �G����ע ųNY '�G8�7;�X&(i�Z}�^�M��Ǥ�ʙ���9�����ɴM�u�$��<�:z�"9l�mw���"6��%F�X�[,�u2�`��efk��lRi�"�h[�c��L��q��k����7����H���9Y!�a����I�|� [�9t���t����Oy�D���xF� �������$vlԿ�%����N%1�K�C����<��<Z����,���������1���D���8<|ړ�wIc��6�{h0�$�m���4g�p9�M2T.g�F���*3�z���3��;r���`qs�YL�c��=�:s��kt8�Ժ�!
� �zs�:�8f���U�-��;N,*�7$��b�̝�����"�N���66u�W+MuAۓ�D�\�����X�V�L�睽�|w|p7L&Z�ׁu��&B��s�ʊ�\Z6��
�G�l-w!?oFV%j�OH����kXF|�ތ푈�g��;G-�#P�+����<����F�6u22�o�P�>%G�dh������w�p'�{�DQ�rP�nH!��%K�crY����&y��1V�era�.u��&4���j���e�h��X�2�H�е��HC.�WM��7Ô6���|����?����\��jH"`�� 0)L]eWPw4��5NL�S.���Z�`�9q���:4�>ڻsOO)��^W�2�_	��#Jc�S0W�{T���ȴH�ɜ6��g���;�uB�0WY��@�L�/�%�h"�<��:��!F�M���9���z|�
�ގ��`��,c�p�����j<y'�<"sfj9q�H����)�#�ɍ�84Ea$�'�S�#��l�S�� ���Y&t���!W5�`��߂�����(��N��zf�Q4����;�$b0l6�W]n���te�~���ϑZ�\&)��y,yW"���P�|��{�1\>��\�f��p�t
���d��&lex_�@5FE��ߺ�E�)R�z�ރ�U�'����?��G�;�% �)���kN�����67������[n]x�I��U���x$���d�Ϩ�e�`��;}���@���H^��B }�wAU?������d��o/�cIh�N	�(����ҵ9D�(����T$g,2A��FJ�?��
=��DΗ�� �<^[,z)谝�˦�^��Qp��mv	��Ь ���L+)B�M��;iw��or��h��C2���<=�o�d�}�Z��`}�Uc�+��0&��Q��������ٿ��YS圣b��P�Q����q����h��~ad�=M�Vp�����6U�� A�7�)1���բ��[J/��[��e���柉�`$�׎����LH�Mmb�|�4S�)_�V��'܊ l.�ϳ��U�m^�T�/�uEh���KQ��nhRn�侇[�:g������?�\��������<��R0 �3 �1�d�(L<=�^'E��ƝT}��4�{�Vgè��|:U�l��E1���������4����2ފ�/'���|Z�~t�M�Ff�I�އ���p+��R�y���Yc�R����tcְ�'A�-�����Z]�{��A?7�ce->��u&�����Ȯ0'��u����(�P>���E�����6����-ܱ�]>5���,S���g����[xf!���Jm	�H��&&9Md<���ܘhQ� EdB~�����P�c�H�T�fS?�Xݥ�qH3�P�@��[,%F�Tt����iy�A{c��j�	f�`	ʴ|m�I䞾�)�����u�c/r�G+�|}#!��aH���v"��=��� qk}J���$h�>Ԝ˸-��
㗓��s����� I��é;k���WOrr�ҍ��Dc�D|�ɦ�����4�M,� kt�T"�,�}6� ����/�j;g��e��TH(�v���ad.��::���M�k
��'2��5Z�HT���4p���L�k�� ��ɺ�뽨���H�D���7�K�3*$�K��k;��Z�