��/  ���yN��	�I΋o��l䢲CwJy�wL�Ɇv ��I��A3N���S�M� �;��h��|P_�ҵ�`����׿]I_���sO�॔�:�\
�w��}��M���=���or�(�be?�42�,�ɵ�m� �>®�$Bt@FP<���~i�q�ҟ^��<�J	9�yI۴�:Sހ?�!��mbH3.��^;�b1�A��Y�Ǹڢ�n��0-��$I-|2-uq��{���E���$��/�≦(5t���N`�W�jddl���Ҳ4�ň}��׫/`;�Q���8��.��c���������#�"O�b������0*z�a�.��2��:̋��iV��4�)u	����\z�1��ހ�R]�/ɕa z��,W��T�X���\��{I��Qc%�"�>]ZG[�"�&.��xق��=�U����9�@��~�u�/Y�l�1v�~���}�ƭ)�!o4��	xm���B����nD\��]�w�`"�,���7��dAb��dm0�9������kŠ�vEWv�C�aa�';�c�R���e,���P����:E�	wz��M���6K�3�]~)׵B���p�w���z�E�Vl@��+�<?1'0b���o��⣘�2>o%�rTk@�Q3jH�e�UV�VKq�����y1 T\�����(8SYDov����3)�=c0fgl_+����/3�0��d�s=.)PJ�PtG�w�l�J����Ә� en� �P��EVle��&��C?/1@������\yl"n��T~uʶ����%�ft������nV��?$�z)#�y�R�~>4�b�-y~�P��}Ǣ������玁����f���J�,����)o^I����Ϳ�~�B5]��K�r�6�*�ƅ��=gP�f�X~'��Sn�l���<�ؖ���������4�Q��vG�,�����5��T6�ڡl���R$�ڽ����:����MހOd�v[n)[\	� -S)�}��O�5P@�
�U��*�}�k"�+��_'����� &"��s��ET�u�_�'�$��<����Y����$oXj1��{ϭ©̅�1��)�/���!+������6���'�U�Ka��p�o�{q�\0�ɔ�*���0�э9�%����)���o��p����5%�R�yeL��ܢ��tY�Z{��߹�>Av$Yu�p{Ym�z�L�o�$.'/<��-�}�]Q6����+�5i��ߥM7kD��rQ�O�Hz��Z�e�	�Vs-`(R�R4�T�/�[n�������l�|��4�.瓦'��*�T�*
��V���k7ۂ1T*2�������N�m	�/Y�H���=
΁)Ϡ=mՕvђ��dp�Ξ�n+: P!��r:諁�E�����@$U9 �Xu8�)�[���e�{�'���D�指N%,YU�T�FA ��b���G7�Va�au�g	g7l�A�������r�<�g~������`ȼ��d�?��"b��1[�D�vA��l�w%A��+9�h	�~�φ��| ����dtl��ݍ�y�8�gp�=8���;9�/�	�$���)δ�I �2�ru��*1_�J!�%�pV��T�0��HV	�<�,�#��}_��7�-����c2e=A6Se��-���B�t�L�<�qh����v����-�����i\:�e�u?p+�� *$+Eu�� N��RP֕�1S�Q�F@������Z�Z*r�e�q�.�}M>܇�sr��爫Ֆ	{ѝPP�\��q���
�[�yBcj���)�guU�;������������RJ	x�׀O7��"]d�	'��9����C�,��lq !w� m��\I�G�ȵf@"{��AO|WW��,��s�;��3&w���R&c�JD,?�x	�Wג۸?�(�6�I���{��s��7
�:�p ��6�\ܰ��֨��� ����%ϐ�����-N�ܬr��v�|LP�l��q�m'C�\"�X������d�)n��W����&����E�"���Vٞ!�;�A�,E��L�QO�����pU�uL|,n���{�)����G�T�A�0��Cr�MdA�:"���P!����&u��Ʒ:��p����O�U����p3���!�R�T��JZY�]z��8N�.�A�i��ؚW����VFQ�&�`�C��/*D�v��T��X�7��)%�{�g�8&\�7D����-9Y�՞~����3�0�]O�w����}9��4���9��F�\�zr�l���CO?��
���x���נ1�c��$h?����}��n�����7����0�*�����lES��m/��x��&�De�&��
җg�7��֞�J���SE�����N�e�{�4�g���n\�'��V���@���@͉����7�邛��b��.[ބ�<�E��q@�K��;�8�f��1fl'f�/�5���\f�
��1�?kidV����ٴ�#��P���Ec�~��j`�+� ��t�S��C��B�g���)��q\�wxT�c@��4�BTA4;�l}Ɏ~K?���Y!�v>������6�"�SƁj$F�0f18�BW��N�����Z�����qpx�c\�6�.|�w�Y(�̯�=�|6���0]�Q6	��p�|O�����.@�i�}ʧ�d�ev����ʈ?0�7���n\Q)}\��O<�����#��S��Z!�9�m�0\@Vc��G>SG|��m4���7����r�m��C�d��K+�װ����zw��GX������Z�*�B����+~�G���>@��	,�IkY�3�TY%-7޳d����N{&���0��u>#�&�� ݓ"���̼��[ܣ+�4]-~��(��C�xOnX�4r�������#�`�Z�>�9ͱpq��F���@m��26J%F��Avn[h &�h��xԙ�8R�����Q�1荒��V�M0�(�|&NH�SD\�G�R0ĞU�NVtr��}:��cM����&�ש6-�ܪ=��{pټ�A��to`�E�p~x�a<���o�2����:t�W���Z��]����X��q���10�d�+�}I�z�N���bkPK��#�������_�A�>m:��s�Bl�ە�ݩ���USK�h6�S2�����YC��m*1�����ޘ8���������"�2����L���t�IW� ���(�YNNۛU͞��������(N���±����+��m�O���D�IA��ӷr��v�N���u)j�.���d=��#�㪜^� ~Cd���=�w�n0�KI���:���7I�Ա��j^*���QԕF1��r��0��q, 1v�U8X/Y��<�hp8�t�/{��w��7aB�0~����8�F�P��'��	�?������o�(������Rwl�vxm?4)sqA�����#"cYĶvŒ�$�BYQ�ɕ�m�ZV��Fѥ+�ᅨi����4��A���_��3xع1U~�8R?T�� ��9�6��'K���^=>�2���J�1��f��U��MV�s�յ������ok�j�w�gc��
*?�ģ%g��{���@��)��,Ҫf�a&�T��`����U?J�a/�|�e��6�Ev`~�,�%-�<��M����������r��N��C�c�B(��z�Ȕi�Cԧ(��vMi�?�'��[���ll�7��0[�O��_
M;`�%l��}i[(����UVӫ#�VuX nl����c�(��h~�"��;U�b��00��*�g���5Z�!�q�M��X�k�����XB��d�A�/�k��n��Z�Rh�_a�9���2�F�����`��g �t��+���i�Q=�D�ٌ�y��~��_�9<z�8u�m���*����gA�:����9v1p �۴�Q��:�����?ݸ�?�����·Gf6��4q����fl�G5E�8�n�7��E��6{�d9�[�%y�,3$Z������fH?=FDth�@��Wv��!�_󧒰��J��٦Y\������Qe������Ԑ�6�;�3�7�q%	�ў� B`��s=')0����$rԑ��d��[�A�����#��+9��`3�-ho�D�S�^{58<�[���e��G�o<H�O�`�$��֒��:�Ch��~��/�x!cRΨ���X�;sIu��!��3���3���*���'	���e� X�o5y	6��z�V�Գ�����+���:� �R�4&ᾁx�>��4�pgP͜�t��'�W�z>}ϨE���R�3����F]X�\����n&	�� �����M�u��!3�7Oi�E��e0�_����o�Ob
��-àYڢ[��'¸���;�lf�₅i�GD�A�m(2�
���r'��*�hb��G���#�0��9X=���#9����k�P�T��"�D�!a�x�y����E���Р}�%�&�B4W��[�����#ŽRS �#]��N�!����ebF��F}����U�Ĳ�[և��h,�H����1ΰ�YZ&�gRk��	?C�s�� �]�]G� %�q-�}}|A�=u3
���nmV��_�����_R쓱m�c��F֐��!*�J2�ǩ�Ӂ����@ъ�i��U��<��+�Jor����h��r�d��ո�m[	��+h�Н9�܎3I�A���@�r.0�z8�~��.�:��`��,9�n�%�iKu�#�06�>�	SK1�V�53���MM2;�O/��"�Ǩ֎M���z��5���N��N�����x)
~l����OE �]�N�~7L�`NPT�{L\N��ɀhaB>�E1�[+��Wmo�� ��/߭{�����F��4#g���⌅���I��� �̀|b�|�{��i�9A'��u&�~�G󦡆f�k��`9��"ø�7�d�'��'v�����U�BV�0y���8�W�GÏ����ZL�O�IV@k�<qLdD��&�6�\ϳ��%;V�W��+�j'm��h^�K�"��?�*�w�-�~F���
{�b���)z�/����I�oM2���l�FfȧZ�u��:#�1v��XY�v%���&�(<Ԓ�qr_��XY�"��ְs	`��
r�!��&��R(S�ߔ��l3�k޺&g��Q�MbF�!61<����B�!�F(�oh1�U��	��U����<�C����8WS��g������Ź��`��x+��4�D�eK5~�!�B�Ol��% J����C���N��i�G98Z"�{'��Q�0M>�t�׆م���J����^MIK ��i��V�8�%�s��v?��߃�	/�=?uG&�nK������18�	�;�XLȁ,ư���+�7�Gӱ��Ln����Cb"�]@0C�����0"�8/A���2��*��F�M5q�Kf3^O0xU���9#FD�a�>/A�6�&e��y~UR �ђw��$��X޳���W�tU�yg�h'�^���Kq�����)Dn�EK��n�,g�L �B7
���a��,�6`%���P��yQ~Ĉ�u5�B^:�����J��& �}X�\����k���-��0�=7�z�W����9��Hßu@<�b�c��&a)@R��ф��s	���k~n��i��%<6X#ꡬAJ�,�E��{[�<�#�A쿥��r�gΝ�ޛ����!��W�_(2���wZ0��v��ڡ�Bٺ�o��[��!�"�%I�ݛ�����3.�@9�M�#['���(�N�.�G5E�z7�o^���\|ݯ�p���X�T0^>+G �F��b�'�]�����j�C�Ur��H9��z��Me'�j�`���EJ���w�"��JCY�3���J����5>���{$g��I���IKRؖN��!RZ������4�E�E�V���Ȃ��߭� ��&t�7u/[����H�^��	+gk������U�N��:���)�9�