��/  vp{,���q�����}q��A��|����He@L��W)Ǌـ�v2��D��Y�4'�?�_Ԯ&���>��kӧ�Ih��ߣB��vC��；��� ��l�C�AIK1Q�k���L+1�J�%I���}<~��K@t� ��r�I��y;�a��x��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<e�2��qK����ﾽ?�w3�d�,�5ن�Ut�"�~G?#�����f6�o��tݚ���3��5$]Xd�m�ү�U�|cY� �Bq��)Cm���;���sU�����*���9�ʇ�q�ǒ������XPu�c�a�����w���_/�����PLf�M�_�	犟I�7/�3�Ȏ��i�~]E��� ��}�C�b$a;���ʲ2�A��"�I	Ci�	�ųG:��r?���~���(��>$mDS��?ã���O@���*��L��p�0�'j��b���K���K.ᵌ<��a!�Q�\G�tN� ����~��Tjk���u�ț�������.QM劻(�Ф�n���a��^��h:�R����v��,�m�y�>���>^���񣙄_�e��l���XMӝ۸׺wF�	�-�����?��[�z�-8$O<�>#����"���hE+�+������\�d�p�$�/ۏ����|���ٺ��Y�+��F�h�qS�O����5>���f��V�j1I���l�C��=�� ?Z�2Y�yr�`5-�?���_.��5�y���^{Z�d���ׅ6Z�E��&ӂV-�����>o�e�i�g<P�X�eΉ!�M'�3gŢݥrQ�e���Q4��tHhNj�R?dEĽ��)���R��A��ë� Tw�P�<�5K���K9N��8�W~Ѝ}g��q��ry�q]��H��Nu���E���Qۇ������}���ܮ�h>�_�v��g�Ǚ{	�1�Z��h�I2�[��g H��x�ݺ< =-'�j�	t��)@Q>9�q��^p=<��� Ql��4?0i�<�`��)�U|
�~������S�	����Pi^�ǰ��3 ���c����p����e��rR���>sH|����pų�V�g>2"�oX��J]<�MNb<&�KTc�b��Y9G����kR,L���z�#�V��	�1��� ���ctd�#��r�s>ރ�ˤ{e[l`�SI�T�:��٢�4c:E�a(-�nT�/$FWR�q��o�`�����R�o�O��I���D �fGF!��ʥ��}r�z@�~�FH���Gf/�LU�"E�ꆡ�N�=�e�'�ÄOd�&V�Y,oyw�1�*��;Ն�����^�������艝��XS�����rF&�ߚH���V��\\��<���6oe��
�^��i���E�-��I ��-�
�U���"�^T��w�|;���}kf�}-A�NїE����0�ss��W��Y��f u�4r@���
��� u)f���<��M)�63��GE��ضSmjp�ޒ�FC2+_E9�nD��h��+�X��C��;��ÜJ�H���Y�Y���o�9�������-��;t#'��Ow�׎���z�d���7]�4,��R6��*nX�:&��%S��G�mT��"u�U�%�R>��Il�7L�g����
�������A����T���sW��mKM�#�
�{1�x�JX��a��`����2M5˃�H�R��:��]0�,р3`��_FK��pl�r�����	Rm	�'���_(�'�3��E) ���+������E�&��	�N�ÕFk�ȳ�<�W ��?A�1���*g�0���q���'tn�O-���>%��I��L�3�qj���'n�m{��Q�0���*�����X���N�{V�����~�,魵�k�Y�>�d��� �5,7`����g�(�M�:��*�]\��E�n�3:R��m���l@)�����l��r�/?�i���Փ�7��{�>���`t��w�OrQ'`N-�	�^!h�X�R��6�����%iJ� ��˹��Ϣ���sp�m����E�F�PT.PEM��^�*F���ӫ�{��� މeP<C���.�{���ѭb��{@��q���ab���������vK�Yѐ0�Z��J��S����`.�x�A~�A�i�ٔ��(n�S��J�����u�,��:��G�B�e�4~����P�'�Y�B��N��wī�0���V�MI>�S�v�. Cv����y�| �����;��qs��N�����0G�:h���+c����H����g"�++2ܝ�	�Z>����q�yeįZ�*;�ɭ$ꃮy4��L�J$�G��&T��9-�b�Uih����>*x��w�'���/&��Y�+��^�1�@'�h���'pP�J�Ә����&!7�:k�_h���V�6���I��I� �p\xh��z��%�_}D�P^W�	��=���a�o\b��� 2�Q��W��Uuk��D1<���ۖbqN���ɽ��z�!qi��+��1��|�{�Z�}%�} h_�H�k���H �����6��?k���b؂�Ɓw(��#	;w���Ā�y]z��9�FQe�R#�.��Wނ+:�*M�����1��E��49����B��� Be���f��c�.��{~G�^�"9.u�-������[�^���{�yT%�djIDTZ���o�[H)�;N�œa�c�S_o��J� D:*��\�(3m�z�>��&=G��m��W7}�2Z /j��7l���c�,���2��a���j�Q��̩��y�L���\=�5 �CVU��k�5���HA��|Z��#���Ϲ��Eaa�b u����r�k�(a�@m�V�S8wq2���c��O�5#Q'�@;uN���b��q�N��>�-�%����T-u6��j����,���9��w�o���#b�}���Sp�{¯;7)���YYR(�؏�-K{��!*ڙ���F`C|��]�fۜ��c��No��Eg2�������+a�6I/�c�"R�Fok��U�N�
��,ȸ@��[��K�i.<��=\hJ�K	���xX5o�U9d����A~ObG��o�� ���ɓX� �x�D��3q�fJyD��B����'��{��N7t��_=�B���3y�@y�-��x-j�Pa��m���y<����?��ݕٓ#���a�G�����Yvi��(��
g��z#KS���h��b�1�,�쫳�� �"�N(ަ��� ���?un�t�P�G�� � ��[R���J*,�9�uY�tU�\�y��G�kBu�D�K>�V��`mdR)��ͦ�@��|��>��Dl����	�OG����VG&?nKhj�8�ι��(+)0�IBtp���� �*Vt.u��.�}
c��,d��ԗ0S��Td��s�sM4����4f����;��"��]u�c��P����\`��A?���tْ�s�mSc򞑡�%7я��~O�����k~��c
�c�\�I�L�.��}>��D,�L%�э�p�Ƨ��([ߝE�I���Th��1�2���"<��3�>E8�X0yB�#cJ;�+?qa�z.C.ɩ�X\������L����lPd�v��'X�
�������K�2Z���Y;NBx*�(7�Tn�a[���MX��D+y����g���ט�z�O4b<�p�'~z��Z�m��LZ�b6H����_lĿb�B&�pv��V�Ǆ�$j��O6��SorvNå.^�,޶�q�k6J�!��O���ņA�P���uj�I�a���6=���K���&e��DN�v-������5*ZK�����U�0���1�[�U�_#mRt�G{�
vĐ��0��-9[�����3�CR�ە�cqs���1��)1+ΐ�R�(�p��*XLi0��OS��q�m5���OX'�ӯ�U����$�Z{Zw~��N�����f2�YJn��Cp;�h� ��F$`l�+�/�3t)>�m��o�N��.�z����@���o���%���r�N}}ߤ��<~N6_�t =w�~?�����#3$g���;�d�a���^�����s�t�}ԙ����ț{��ָ����B�zh�Nŀ���Nf>+�����Y��2��j;|l&�w�}VH�������ےh&��{�t00/��]+|��ꕌ�K���K
�G�R�Ȩ\��e��o��4ZW.�-.�������hg�D��id�lt���}� 0�~�03|� I�>�@F�hg��c��	�h�p@+H�Y��=uUS�������X.��j�����ɕ�d���Ȃ��?���J���)9�zV�����:.O�?T�] ��x�W�m��LրSz ��	��z"�Ij.��}��/֫�.��$�%_�B$w�:����Z�օ��eƛ��\LS��0���ok��rK�&U懖��&��p���Qd�
�+6��t�X2���L��
C1���n皗������M���W�m.��l��2�e�0ɣ���n����F>�����o�M�k�?�w#��}9j`q��U*{�9��!(��m�K�(ߵs �}���� �����G�"}XH�ӝ1�'8�W��1���F�]�j���vH�!3+?t��,a^��EF��@��l��e:�'i�L�s���O���]��-��x&�B��q��-3�r�V��t��t�v&7���:����2?�(_.,�2ac� �to���|�uI��X��<A��Pjq�h$QN.&v�� ���{����*�z�X%_�����s�| �v������jG����`���g�����j@(2���z�%J(~��jr�Hz�i���{bU�в�:���-qrT%7����X�	�����{]�`k��V��.��弳r(�^`�� �σ�`��M�(u�LkuD��ʚ������{�N2����@�{���7"��c��<dچ�kܷ"Ĝ�����MGH��o�`=���>g�1S��,j��=����05����}s��d�|���H����u�l�<L9[���D�O2[9��l�}�YJ�F6z>6]=N�J���5(Ð?� ������O.���m?��R(1 Nz�'��u**��V�E�q���c<1�CT�d�Q�����=A��.sù�]\�C�]�̀	�;׻7��A�������~g�Pq�Y�0�ɂ�xxO� Ar1\�&IZ���T���BH��[���8{�b�&��kH��@ڍi��Cʰ�>ԪpA!�5��zNꨎ����ޥ_tN�i}�b�\б�fbU�����g(\����S�`���܏�'c��������m2̮ґ�L���(
�R;�<���'�k?�>V�Y<�@yl�,��Tj80��v�P����~ԡ������b9N�v0&�����qNZ�Xs�ő��BK>��$�"��gVn[']]P��>��H�^�|���D�]�S����m�>mc��������������%T3�����<�TG�Ġ&�DO*��_��G�!b�q�v�8��8I�>6+0Y+��|]/S�qN�T�ܲ|��`��]�B��v�I4�#����LBl�u�/e�傢�l��ы"�]�LP�p����$�#��|���'��F4�Q�νmkjׇ�/�߮E���!��S�=/��󠤸u�����m��0ܳ����s�Ioc���wF-?d�Gȥ�������y4[ĊHwŦ�@�~֌Bg�#�}X�.V]�Z-��a�%fKǎr̓���@��w+g�6�b��%��j>�r���m���sSK��E)a����'ŶZi;�B=�mE�$�t&� ���q�Rp#�J)��W�d��-��DՀ_����ɍUkGU�1_fw3W7+��L�U��	����^���gb���g�WzX��iLp @�	q��z���%���|Y���n`���G�-5S��B`���{���d(i���_j�r�M²`p��p�j�v��ܪ3L�Z	"��
��ů���c�dB�N�]�G�zPԕr>���ռ��!�Iٔ`��ҰN�F�Z+������cǶ0�/�#����neh�����dDe�4������N6q�~P}9��<��A��"�'��
���ͨO{vxB�d����M|�MsI�lf�N��Z�A�*7gбa�) v���2��H=�f������<8��n?"�M�
�3�xJ�����ʬϾDb�0�ӽ�Eu��vfwS�C��R���y�G�9�(�,�[��?tA��Z�k�w��L�k*��a���}CJ�A׈�&6����Ob��[NM��-1Z�2���CI�SX`�7��w�Ì��o���� sz_�[�c>(V0�b����As�@�/J�|���T�i�K������ՑD��ҋh����9�`�}��a� ���2�S.�1	G9xC�m���A��A��2�4o�=��=A�kD��
 \��(Kt&,��������>�Do���զs�#����qL5��$Ģ���WwUl�/����	��>,\������1���[�:X��͟�̬�'U�u��ʹ��0�j+�(��s�Ű�9@u��V�ީMR R���c�bwsmEA�L�>��+����e����{�%6�	��O8��d;|W�e։<%����G.�m)���T,J���&�+�zƂX����X���Q{0�r�1��7e���6<���U�zRm��w}���Z}����pI��L�/�Y��%B�w,�߁@!�;��|td��4��G��������fc%yQUy\�[�q�Cc[,P��(�Sd�)#&��~஺ǧeU��g�u�M|��k�����XA6�g� ��_���K$i��ZZs��q�H�[U���rrm�Pi�k/��u���^T��ZN�X�kw���|�/{j�3Ip�����r�^�_#o������G���(">p0ޫd`��Ӽȹ�(Z��iEj�u�7s�:Z�F-�f2��HZ���w?K�L�qg�?BʱU��I�Y
�ԨH�ðT������G�u8��GݹH�bWxCe)�w����W��8�J=�IgRQ{�����J!�HA�72����3:Mj�T2QK�(��"��.>\i]¡�-;��D"�%���_: $��[G����*ʞ4��c��`c���V�7�#��c��^�]�(ϱvf��{�i{����Ҡ��O�~/�~�#��A�ǆ4����;3j�,�~��̌�@X�È*k,g���&�U��SD	�5��KrA�
*$4�f�o3�7��}�>L>V�)� %!Y�O�8 s����D�T�bs0������Zl��Jw��d�˞"�^��)3���0�r�3B��3���t)���2�R8�F����2��7-)Q���?4���8��"`�`��I"����؃��?z�T#��(ۄ�tH���7lp��]1�����^9�L�.Ќ]����J�:6,��	�<�������B�p�T���������C��J��W�G+Ӧ ���"�*�n�<'�_>�[˸���J~ Dbϰ4凣�^���QɊG+��y\ G�D4^����%`zq�WHq?���"l	���0�Ə��(�.	�%ȋqds�J��A���:YX|k�'E,^���h��B�_��a���ݡ t�,-�#������=	2�B�U�\�8үxa"�����$./���r���N��x�-@5Z
�'������~7bs���X�����E�V~o���7�.yFk��է�p���3�!8�8��c�E+�/�'\<o��@���s��y�⹡<�𙿕t�һi�.k�d_ߓ��9 sIF��>l��-�t�n�x���p&J������za���oH`��@���P����5�"�5��ܾ.������x$��D�ֶ�XF#=q���q���Y�$��R�TS#�=x!
�6��q
�B�5)���#}�V��BU������<�is�@<��)�2��u�4Y��8��ʆ�J�ں�� [=ۓx��ȏ�O}:�!�\�n��X�Z���Qv��a���U�\��i�=�gy�7o����Ns^=�r�شniu�l���9Q@<���(�,[����_d{\;Z�b�3���Hs<�]��&��"�<�4z���&.;��]���}�����wm�	]�2�3��Bȩ��5�o/>JS�Mݢuu�0���������X#,�iOht�z�b�zwI*��k��yL#����0��>�e�yq�(�,r��=i�!��J4l�ݾ�Fi�>J������O,����UM�������\���L���g��ӛ-�F Bվr�u���0�o��W �����g$nW�(r�yMN��|P�I=?�^�a�0��F������W�t�P�0jԢ���Y��#'�Tlw��@�6������S���:���?���n_�B`�f~�'t����$�U�����i��a�.�[[�C��.8�w43'WSp�@�Қ+��
H2�y�b��?"M����4֨�/2�1="@�?�����iZr!�>�t�
Q�P\�1��M�=j��'�El�������h�S,ޚ�8r�3\th��"��%�V��'�?*z��5���8�!��j#�u�/=�0�,��%l�b�)=�.���fā(��N�����ldw'�;Â�]�d����`v�^��X����:�yK'�G���M�T��}lr`I^���Lw+�%_�;���ekᏽ��#3w��f�%ƽު6�ܟ�y�N	�FrF��KP����1嘶G�;`�0P��4U�ʂ�_�_~��ܘ-�߃������lN� �p4�����(cw�ۊ�4��ڪm�W��G�6��ս���d3���_&	��#��d9�����qnň��`&/Z����:U�Y#p{��*5������_��$�PJ�5TV��vDGQ����̮p9��ğA�~~�r��\�/��T�fG���@u��+"ߕ�ϝ�vF8���@���RA}�L��B�:}��y��f��i\y1=��=����Z:��#��G�� ���`�;竂�>�6�!T�p.�KL�����²7�_^I�f-�H\޿�����R����� y���SԔijφh� ���r� �,fg����yngd��Lj��Ɖ���0�5љ��*ay6bW~8Ӫ�|4�����
�E��F��d�Z�����������ͣqc��$ξ���o9��jo�C@��:��d��]�&��G�# 8.X��ך�~!���1�/]�Zjت�<���C��3Q��:�4M��$"���l]�d�� �3��z�,[l�A�Qʢ��m��I ћm ٖFK;�R��5��,��ĻCC��fə������������p�r�`��R�/y��!��&��h�uĸ�[p�6�R��h�<�In���ۮ���}���/R��S���=kF ��on�P�����ih�|�y{|�YQ�o��G��m���s!��&��:y�~"�a�P��΃�ɿqA��QR����F������Dl7.Ct$N@���
A�Lհs�4�[V�M��IK�s@���V!���C����{tUG��K�`Gy���eOPU�<��I$�1%*n�u�Q�
�lI��&A��9̋�|�1�ྯ�d.����E�Yn�)���ia�ˢ.:1�z����^��2��	����ܴ���7W`�Yt@@�zH�^Ǽa�OD����LɗB��񖨹��SP��q�M~_n_�J/ٙ�)��%v���V�I%��e6Y���#p-���y��'�_��<��Fk�v���$�+V���&`���>k<^�4��q*�$����2��q6\p�� v����Ͼ@K4RG x� �sH�K�0Iz�㻗�Gܞ��í:�*P�����X1��l��j�]{W����52���x7�^8R�<O^@���Μ^�������ޡs�
�둑[�Ҷřp���6�f=	�)��\��t��3��וe�L��򰱂8S��eb����ֹ%[Ơm�;�rb���{R���C�|�o��`�94Rj��j�v������o��|��H�D�X�ߤd��h��fԝĲG]�z�c�J9�a�9L3�`-�;G�!��n�O&Z#��̓�pOW��v=L��1�C֋�{��ԟ�!|~�i�.��-,0}�� IT?j���mZ4��2w<����Ƣ�u�ߍ���Pd�`X�n�3� �vv�^bV%�l�B���A�q�$����Ln��D����y�;V�߰7	J��Nyj����\�^ ��h[A����?I��
H�i@_,���l�юj���� �N�[L�z�����g�-K$�jG
���_��c
ꀙi�n��&j�zA]2*��B�O�˘�0>��lU�N��M�@
�`%#��[mw6�>���g.D_&�����W��sNw��ɩ{qZ�X��0��BV@��Xg�tJUWjD,�c�����׈���C�䈑r�)���?��Q��|4h(�_x��Wtp�e�s~�E֡ǜ� zn"�3WXـ �@P=7m�V�gǮ���e�^��Ȩ@��`�u��W���s��ֻ@�U��8��UV�_�E��;�8>	��X<�ͷKfP���0���#G��mp��Ճ���V Zk\�G:<��FkEN)��,��'�Z9:/���W#^�C#�km��䚘x�J��"�[�Y��n�� b[�ch���\N�Ņ��,���Ý��H9�QS_�O�;�oԥ��r"�����&�h^��(�* %>	�Z�Xe���4|�bS�/�Ֆ��Y�2#����C�wdH3�E�Y}�7��d�GY�2+Ɩ��^a���.�F:"�}�M呂1	�`�M�U)�P$����R�mÛ��(�Y�>�c�*��W�)�+n�N���-Nٙ�Y���S�1mч�&�OT����\ �4R�B?
2��d
�ֲ�M]�ө^&. ��?��8��˩6�-.�m��\�	KpvM=}�l��Y%��$h�fECX�(�3#���R�Vy�{�L��)Gjtf�ǳ��3�aɏ"�ƀE��;#�,��IhU?�2�d�3��E�NS�&'���}3��ܗ[����Y��z#�d`�qO�)Ɍ�z�]�����.Zq~f���=�~���9h�ӓ'�^Q>k������
=�!�擠�RE&�����c����z��B�̞ܭtȗ���-,^6�*/QK$@�����5�8R,���p�O/�|o۳���A�Ep�
 �	f��[��05�!��<{'5�+��u��k����2��F��J����۱��	D��c�WS0�D��D,w���B��Y�/���i]'�B���vAH-3h�Ƽ�N�cՄm����q+[��f"Ȣ`-�D��m�܇4Z�Af����@�U>%ٗ�@�uEg�ؽd�~� b����2��2-���܆en9R�Ў�*�����اQ҅�^U�P�i�n�"���Q���|�$�'��(;&
�A����a��\r-�s
": S�I5�r�� ���;h}i�<�T���%�����g�]8�8�~>�D��z�&�������
�̝N�7Bm���h`���H�eʄ�)wԨ�,K�7���hAE�Pm�e��S��(2�%��Sb[���!��`Lg8AcL�a�Nhݏ'���"�$l;�b�/������S���ء��M�C��D:��{q�W_Bv��,�v�z	�~B������*湽������{En��[+{�Ы��O@	�sr蠛r����"O,���x!�/�o�Q�ma��I��w:߉U��4X��v�'n!
��Y���Q��?B@�Р��(L์�Mι�͵h��9�w�z��W�n�FE�3:����'�,NEr����		-�P����2_\�!]ׂ��D5�4�w�9��%s��4I��BG��E���gJ���!i�W)� c�KBd���|�:I����S}��n�W�g�}�t��sc��Ƥ��mGF��us����5�B:[{:_p�XD����U��o�#?%�0S�����-��sF �:І�]F%��^�(6����cͺ	6�"�d��D�#'�3j�O�Y/��,>��b�[G���t������^?�GnK���4�� X̥��Y�Q���B��cF���G|6�'.�4�Q TƓ� �x@�Z�����)�����u�q�'h)��L�po��m�6�i��P/���?��gBK��%�LZ�UX���XGK�J�!�L����3����!@��Q]
D�I�X%�W�oOW�ӈ0�!読�G�r�n��������tޞ<T%2�H|�x��&���e���d|'��O18��t�=�X�]�S `���eW[�`���j��v���<*�d��IC^6H{��W���z1o:r��E}	�F�^k?�h����7�Gl�j�X�������۠]S�w�c�|�i��u�����js6H���l�|2���	x��7q�\�P�*�y��B��v�0/��.�p2�H+�1�I�S5�(2��@����Zx�yЫ !?�K�;����g�Wkf��ƴy�:�kq��t&8
m��I��)���\8y'�uT�Ӏ�ㄞ��&�R�`�S ҅Nz8"X�"���^ԆL�a,��Y��$��ɩ�40!�y:�C���L���cW~�n�ۋ�:�m��~+UY($yq��a�`������܈�����-?l�}]ߍC7)�)�a�5�"�#,{AS��҃�0��uڌ�� j�}���'(�gn�4D�c���j���{��1u����S���2W]ک?��*cԙ���PR���j����� Q�n����l����K�-;ϠY���Q��i��rQ&���Q�=��nP
Bl��æ!6���L�c��#�B�֔�y?漍�¨�}ND���]\@P�_����^����/B4u����L�lYPp�FlI�ݲ�w~��Z�L7�B��>[����N�	FdvX	o��n��ǟa�hR~I,��W�>��ďZܭ��W?�_���(a������U� U-���M4�UfU���)ىQ%L)��U��$�}/�c�?S�˕fvSdLS%9L��5H�\Y��=7�G�ٷ�S�uJ��z�S��.G5y�;�� �L^�.6��ȡ�l�wEK$��s���"�#��n����q���V���]�һ�)��nW#�
�\^)�1�dN�}�������ʱt�X���ߛB�8��#j��Q�+�c��-������I
*�|�f�~#���|��8�p�
�]�����=�0:�Z���DK���"��4(���ֺ���""���^T|�L�!-�ͧQb���ǖ5c~^����|>d	���?�tF�':�dcg��4r:�����<,|�����QCO&���Iq�y�-���D��<��������(���B�~����v���Ȫ"�����b�I=�O��dx{�υ��|�&�~2�b�(�  X��f r�,t��t0��LMN�H��������m���n儾",5�3/����-l����L��|Ђ�5*��u�m�9aMꔒQ�1]�1��T�f�m?��dޤ�Y�/hDq56:�~ת��I�W���߂���y%�E��5؂�|9�&�֣$3�1��6�%&`/Fd�y��N�4������EC4D2`	