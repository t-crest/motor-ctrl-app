��/  ��w`�L��A�C��������W�f39>ጚ(��'�����s�.���9&N#��5����\<
�Z��Q�nZun	�_I��$R2kc��LG|o��;�/�ù��9{�
��'9RW��
��j;:��w�'��(�w���H�������)
>^��<�J���6�����֕��**�4�`74$�xe�#]/,U��C�Z��4�&y�,wlK ���E:�3i#�e���N���i�/!t��� G��Z|�m_�rU�lU�6�  eTpO�م׻�>?(<�Z�f|����j����(��D� �h�$�3��:����zH=>ǝ��+�^$A'۩=��������.φ�M(,�K�OFְ:5H^�~���i�&��+�g�5=��$�w�3�J�x�:y�}�rd�{�g6f�k\7�J`���fD[.¯:��2�gf�N�}�y}/#�Uа�N��v��xq+��q��R{��ܧ�<�,q������E���
��ng��������7��4��Ʀ�wg��l�����?�ޑ���i�k��q	M�}h}����a�O�щ>/�̅�ޭ�җZ^,�fY���_{'C��8��W*����#��\g���';�w׻Y�#d������&E�{,D�j5�oo"�QF����۷��=�|�\�:���b%�i�t`ҋCY�hk��t:zc�{�/'�o~;��ZT�Dd�?�a�`�ӆXnJQ���#�/΁0�n$�)=]%�J�I$���lMJ�[W =��x��8%>K�Px*k��ī�A;B���N�Q85gY�7�0G�}-Z�WS��Y���m	�n�>���`