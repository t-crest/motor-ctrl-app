��/  �ZT ��5�K�Q��l�`O����<�w@��(�C͛$�E.�O_7��	�A,�� ��Н�,����xr'���������i#�9�q��®-z�M��o��sM?�Z��7,7��ѥ����]���Y 7���K�w���/.�Č�Լ�*G\���	�d�E^��<�J���6�����֕������h��3�"3g�Ĭ;�:.���VDvaO��m��,�l|���m�Qht��uw�U�g�9���j՟���L�QTՕ/�P���@��Di��흳�8J^���A�ޏ�wb�,M7}��+8}1��@e��f���v����|�`D]��v�*�sH�t�J;ܶMØ�̃^�je�y���E8���J'�ǣ�nQiVȂ�GТ�xQ�˹�{�|ڛU~���"��T��	D�	Θ���^�3=ɦ��jNg̞�����Oa���"�:v��MhGL���%� S�Sc����u��(����p�E�Kj�~B�K ���my���S ��8n�a������AeX��0���f��ܸV�,��`E�yA��֕��b����DY���~f��4�_����m�(S�u�u�Q�z,�O+��{I!���N2Aaٮ���$���$t�u�[�@q���9��޹�~�:%O<�͍�!�J:�,�6��¿��=�OHY����<�5�._Ѭ������|�ui9�6�zi-v��(�Eu�6�x�5��68���/N뉘�:OL�]���Ų
v�s����Q��p�oSx�^r�]�?��\6��fx�U��ܳ�㾁�n�憬�z��\�
ơ&7�'�V�װ~2q�F{�4������c��f�BM��j�܄ �6��!��9�_�@�0��@��S���d-0��g��5��D�Mj��3t��*��`����OA3F�ʀ��̬��q~��vSm���؁U;��xu�Ь\���Lg�7��r��b���?o�Z�G�Ge�S�)�����-���m?��Z�k1޾EU�l};��cbz�Ƕ!ʈ�4������,Z�wii6���id�Ӄ���p��*��8C��>;.N�;&U��.�w��}gi�3P��C�"�K�4�[<�÷H�u���Z�xۺx�dG�PLj����Z�3�
�=اw�E�J�|���91�S՝���P�w��"��"�AX�4e��/ğ����`��ƍQ2�%����{ �0�ǭr��%$F}�̛�5�%�$�Yh����AZ7���A7<ߗE��������W��4���,+�E�[���yK1S��&�'���CQ=�c�%qx�oU���ܹ�����Ǘb�bFa�ǫ��#�K���M�-[��=V�ﮊT��ҟ)�Rڪ�F��n~n�L���0�$��ƒ&�6�O�U��D�1�D�_.p��qsvei�� ����]�	1��e�]�NIHܛ8DK��ɳ�/�T�>��ݙ8Ը�I)�^:j�&�r9<��6���L������@ԫO?����xե�׆n�p�!�~x��ˢ�1/��m��`q�2�|���i��Bߵ#8���s%ۉճj�^��Y�:���!q/پ��z����m�2�<��Pm�:OZȽ5)*M&pvi��E<�s�QF���vA���K/M�YAѤ��G��D�<F�,R��W�q�B��kH�ְTo��x�|O"�a{`Ȓ�Xb����X
^e���.:�c�}4������U�O�b�Aobz�9���"�/�dIdOk�E�(<��8��^1�n�nb��3[�M�\�qb�m!�EBzl���K�	��.���,���q�H��O�^�s�]6`Q,P���՜�9Me��s��a2�ۈ�*볦8��r^ՙ��a�^ ���sNZ�y��ϋ�<�4�>���;�| 3�ʮF8og�"��5t��=���R�m�$a@>�,�Ʒ��lw���*����<�� MB"yk�gV�&s9B�h=�AhIjJ�Uƀ�JD����[�v��f��O#�5�����S�F��!
�Gx����r
S�K���|��ih_�\Χ<�s�̀�0��&�u��+�nm]���t�ۯ��E�I�1N^u�д������"m�_�"��B���x��L<�7$%XX�tpaGn� �6:���@���a�M�����/#(��W�8x�T����l����/�v�T�b$��c�*���{�ك
�ۯ�������/D���6y���&c�- X�3{&25��6Tڠ[3��	�	��ɔ�
�%���@����a}?(>:kZ���s����X��fD��]����?����ƈ�r7�[˖�s2��Y�^��1�5��n +�k�|����� ����n�����MI�ZMuVJP�o.<��p�w}_��2���4�X�(�F�'hGK�i����K�a8uP���u��Ƌ��\>���?�1�����:�]�>����S�YK �j�������R� �j
�G[�_\9�6%|����=�sQ+c����=��M�F�m6��ߊ���u=$ˀ0!�J�_��I�^��Uݗ��T$K+���j���J���;���U^{�W�F'��_���U_ނ$0Ui�y�Qtn4�oJLg\0�M�2+z�)�Ĳ�qDn&��NW ��F���cC�_�*ک4�G�Vqun�Udڡ;�K6������<�:˺�EKEW��q��	��3M��W9wv�j�K?ٷ�Ȝ�T}J`��@(U�*O�#`��n�z:�!Z����cA�)�˖���DO�1F�筎�}��V��"s?�&���}�H9	��Ŕ����oG�4�=���>%��WKU#ɵ���o�>2�#']�� _.��e�_��tS0M�:��DsMH���#���T��);s��3�Y퇢l�"s����^vjz������y�#mpCk��^E���@���'��ڟ�����?G
a��
��<j�"ʬ|����A��Z�?Q:��,s����.�8y��ų�/�c"�;"����A����_���K;���-J��س%0�Ԃ����.gU-�,��?��Į"�/��>t�:���:�h[{���i�JvHr:���s���#�eg81}�(!t����f�CR��N�$�\^�2ј����n'^.�W=���i�s�BB�� �B�@��)`��D_W:��[3���łB\[��.��;�H�~��.U��D�PGX��Ɉ���ba��͗
������^Ԑ�dnĝd�Ll�v����u��]�ѲG�����&��[-��@�-z��������<q���C��VL���Df�<R���B�+��?8B�ekL���W E'�B˞��)+�l�rpR�U{2D�)i��T�Qψ$���8���+���)��%�]S���(���P8oҜk� �vS���2[��=���DrybW&�3cXП��2�0�3'���t:_5�����̾	�J��P�d�~��3�y��A]Qfa���D�U��17'��ì�,�$<W
�-�	�F��9�A��yN��2�}j+��8���r��-\HkZaF)GJ�j�i+�A���e��ù�¬9��S�	�K��̟���Nk2�_�j���:^�����XM���v;׶F0��u(��R_f�aX��5�`F��E�0�=ǷB���ft0��hy�%�Rs��[�B?5CB6Ib\vY�|༴n��9�J����:��ǥ��4TfT�½w
0
�����Z��@4E���@���!��fN�|�G�
8E��s�Ϭ:��~KF NPkI�|M�8�q�-)P@��o;h;ǽ&�S2%{[Lۙ%w�(%�v��q4I}���x��t.l�x}7K�Z
 ����LT�;w��Pvc������N6�ҫȫ�I��b���Ui�E=V�������H'�巰����e��rb�谾q�J@U�<��Q:�
i��ū�����L��l�(N��9�T�*���6�0p���P��ZZ�$Od�Qm����KXVp�2!+����I�p`gvoh��ޭ�R�C)�D����|5*e�i���5��*�A�D�C��˱�=�.(l���=���*C9� ���������zp���v�<z��P��,iN�%�����s�W�a��ڠ�\�/�3Z7d�O${u�Z
'%��o�I������?j�+V,������<�M�xv����{���E�)�bmu�}�q$$@�g�7���Bʠ��H�%�6|����1&��hm�>ػ��H{8�{4hS��5�iN�gx��E�;M�.����."+�"��I-��)�,�p(�L�̓U�dq_ʥ�<]��O�����.�g�(,V����Ч`�X�T�>�~EҾ��oL?��K�3J�Wq��kV�y2���R�ڤ��#�/����a��A��$�B�*����n'�C���(H�uY�V�~꟦�fk��n[�ꉭ�p������I������"�pj˯������[���.5�I�?�oɅ_�l�
Xخ��d��r���Qb	�uo�q����=i���=�0�&��� �9FJ�ˉ�SL�;��K�c�<��\��=^��Ӎ���i��XJf�;c�cE�5g���X��P����.��;a���䆷*%Om�e��إ�Ք�?�IXq�PL��E/��ͨ=\�z���Pf��K۪[�x�@�#�$H,��Fl��d����V�%���<z���/�n�paj�`�����tĶۗU����Cy{'|r�o�x^�)b�ڧx�d�
j��E���;�y��<2���4����g)4Ք��s���������R�JFA��m��}U}PL��F�G��x�U��&��L��3��,��#AwIe�9�!Ćf�m|�MC�|i.��zB/���T��a�ο:�a�3=�3$���B���9Ҁ�[:m��>P�ݒ�Lg)0~�@�\W{3���h'��U�|������ ~;��7X.��l�SR5��9��|	wWS���{
@�_�%7J��b���$
���N��ӷ	j�t'=��<p�����VCV�f�l?�w��ۙԡ{m��b,kpf����N�U7JUVՠ Q��൴�Ib�&	P�cKc�[�Qy!w���;���j?�%����r�ؓ�fl���ZJ��QbEFj���j�󧯫T��H��td��k�mx�O�[���kԐ�:MeŖuVSͨ�׳=*ج�m�K�z����bX��2����)�C�/�P����w��ӏ�wa
%� b3�̈́�Rp������A�O�
�//���9�*�ǅ�Ա�H5�g߰I�jZ�*D�edW�9��#dCF��C��CY�������Z6>����d`m�s]_�\�U���N?N�Y����T���h=~�����"���)��z��Rr�9z��uh���3.<}_��q�pp��ɑ;~���;Wr��Sh�Aҗ�i�E�K�����h�ޠҺ�z����#jRO1ЃS��Hkn�͍YN��ʉ��q�V���r�8ǅw�\ݮ!��2�׍g�6V����*��r#X:��Թ8���|dG0Sn*��/s��!�?��T�)�>��v���#��SC���g��L�1��Ñ�����������l�U{p�� j�'�%��R?�s\*r�& ?b3�<�3��d�#�v�m���8A*�Km������
���Z��&TCU�FR�\Ch��g�Lj��%���1��S~� b��T�/�;���X��y�<��z�Hb�3����M�z�:
���*Z������S�kA׆�>ԾR��b��=O�0��:���]���@���)}�7�^5���/��2i�i��DC�OM����ٰ��: 	ib�����+k,�'^�I*h*^/_��o�|�p���~(�	����/w�%�.w(;ݶ��Ę���4���LT�#J�U���OzhG4-d��/��3D���\Mt�	GiD�K�.i���P���J�tBr��\F��_C;5�I�wc�;Yt�)���G݃������Rs�gRF�����61'� ��nv3��րsNe�3�Ij8";Q�����j�+*����g�t���TΎ|r;2w1nn���\O�SqD渝��gd��F������W������?�s��>Ʒq�͜{���;�(yU-�)Y���Cp\���U�޲i����KD1�/�#�Jg$0�5���:�ͻ(�k��uy�����"/��0M�3i���钤�A`��<;�]&^��Bޖ��P"Cܻ���/��6��J��ۂ��������P:�ۢ�	`�N�d��VA�S�!wZ�'�գ����4Nn5�AD�Bn��:��dwha����I���G����u�mm��9UF�l�Eu�gǚ�!�O�8��>��@�Q5����E���Åï��@{��=s���͍�x;{�|�����@wW�*�P�a1p�8u�3��������;"C�O� |NrA��kl	/V���^a�]��� ���dcE�l]Zd!�k�J����b6и4�\�i~��cJi�\��Q\34�VXT}֫�w�Sf3��	��HQ
d��~�i���>a�cZ��E"�P�'_ŵ���^��2�
�����cyZ��5�͹N��=U����_i�&��/�$����1�)�ʼ�$^�Rnj�ы��������(}�0����/�5m#�&	��C�c�4cR���Yi��@B)vN܄��$A����:4'��wQ�/'����F��q�DK��Ǭ��I������b��&��O8���\C! �6�x�#fM��ts����`M����TMFP�~��`S����M1����>��X_.d�M�/��J	�=�L���|��r�ua�?�d=�����iҼ	�W��K�v��_v�b� �qKMz{`O=uG-��}ٓEO�W��PzL���Q�2%[HR�Jy�ŀ^�(�
�B
��6��;�u��Q��:�Ix��%.���.��^�rZI��הb�I���a&�MqN�f_by��|ǡ�e�8����zc�2�f�t!v�wGc7:�$�9�5����x���o�UUnZ�e;f���Ԯ��齁���7s�*:��D7U�s�1��H$5\��<ڃe�Gɍ�S]��i��ˁ�$Z��g�P��m(L���f�
��������1�e�������TE�yi�Cڡ��%m\S��J����V�c[���z�{�n�y���lnn��Ѥ��A\�8՚O�C��Ț%��0�F�����Zv���7g}����:�����&�������n�()�J����f���=�<T�Zu:kw��J��3[6����`3��e$È��gXi�
@�&%����Y��`ϤP;�M]�.�/�ŧ��\�,����ڷ�8�.(�9�*�n1������G@v�*)$���̋����8�b��T�Q�OӨ�����곌k0���=s�?c_9��K�Э$��h�b�$J�!�5�{��7JT�`a���j��W\å�.���64>�@�xx�S@s�%��Gb�w�Y��@�J3���+��#2�Mt�w�J�.Y;�<.�K�����sؔ�}'�RT��IIAudxr��Tq!�(Z��y��2i�����g�j�ߖcj}�;������9��9 �]p}�G�+F��gi�Pu���xm�=�_L:���������Ҫ��J{�I�M�۲��� �W��1Hl��q$N�Fc*��=�� ��@>ZQ�>��ʐ'Y}$���%�C�S{����8�dL�ddB-�X-|@ft�@WNl�vt%�%�X��AۚV�K��"�X���J���p��,�������Z�a�ܱr��m︰<�G34,1�h�nO<��A�� B�9ïO��νq��Ւ��*�L���QC���B��c�=����}���B���d]�Y��T���CEvl!�17��:�EVz�
��AR%����k֫1�la���KK^I�y�񤡀����C�lzJ��˽�J��.M#��ߥ�F0�(oz��'�b�@v�_���/X�{����U��%Y9cv�C��=�S2c��C!���H��b:KS"����(�Yg��:��5z��Ӂ��2��?��P�rB��@_����$����vK �`(�J��b��k;��\� &B�G�N%e��µ���HI1�4�i�̠I��Qwf]I_|N�C����Oo���S����#w���lk�#�\pp����j�^�ϴ�&(�_Eǵ@��m&w��/�F{�zGqh�Ē�w�Ƙ������Ý ����h(�G^�SOe�Y�q����[���P]���$�F�zy2ǫ�˻�H�Xx��-W0z�C�w�ؼޡ�]V�8��W��9��`>�h�ٹԎ�^g��s@-�U��+n�r#��B��A�)>2zғO���A���^��U�D:��p�csSiWwn~J*��K������ɵ*`����;qkk(k����#�P�Ѝ1P�.9�0q5e��][�vF�zH����[u̣_.���v(p,A���xW_?M1\G՘lJ�|N�<�=�Ҽ���1�+���b�gx�:�] Aj��[;c#���h��Չ���w��Yr��2/���hj����� x�zE��x��й�A���D"SkK��ӽf{�9�f�:�t��e� �i�~Y����-�i�2$"a���b�7��#A�<��v�
穘iUNIa��&OH0�!ĪV��UY\���0d'�b�1L)��C����lor�3��y�=_p8��LyU�rS�����s��dʔoPj�5�tm;����˃:$+,8�l��<a�Kah�X���H#b#~8E����Q�bf�)�l�g�!���N@���r7l���L�Z=M:����7z6;d���C���D���B_�v�ӫ�G�:?����ucl�0VM���ӝ
U�W�($��@9�^�X�RT�a������n`���o���.��S<s�Z�Yc.�f�֊��x�,���'�N��l�px������Y�F����gW�xMb๼~�g?�Auf�5 ���"8w$)��n��os�w��ᢖ�ء�ˤ^�jv�	�r��e��H�83rj}x^�<���H��n�I[8N5B)�i�i��5[�+}�o=he2ºx0MQ~��b�(��� a!�$P���Cڝ�G9��U�� �Tn��C%z��`�o����ښ� j������5M�! Ox()5��ܒ�Υ��&�A�P14G�;��VxtH^{0ۃ=j��\���p����x�������U徥x�f\��m4nh��T�#�o��0Ip�~�]B|g5m	f��N/&���	9�&���o���n �����Y�4�{���h�\K��B!)��>���`�:Z�JȦ�i�?�[fS��!���Rj���@E��LzD�5���G��qZ���$��mc~��)ƀ��9��L�
��G��I5x�O�R����B_�[�&I��>�B��^^�զ2�<��.��Ϝ���%���@0I�!�uW�Ig�)`ԕ�R�VmOM��lZ8+�Ҏg-�j����^�p�kf�-ǋ~d�CN�؄�/�c^�������!��K�����V'�qUw���a��&��&J�]���"���5��y���+�t�����=���T�|pT5gv�RO9i!�;��$m������kr݊�L��`�׳Wv�!���	��M�WѺ�X�*�T��	`ԔwĵM魴>t_�D�L��p�9R�ƿ6��OQ�M���-�ַ�!�n� �Nn�{� $�O����>��ks�P�^h�S�� ���{�J�7�	��](����\`A���2mZ��&�^��7Ծ|fL���@��Ǥx��@��8��I�����ࠅ��n>w6���\�M����|�v�P�� E�`�P9W�t�eV���9*l�z����U� �'o��&0����慅i��./�3��54�A~�Z�N+����Q�L~��N���JN�l����
�#���+M�"�Hs���p�c�n��*�ZC�	�;�����k�~��0h2�UO�7;zê�����,����V�>�2�8����ҵ�����([��#|�4�9��U�򭫾��嘊j����*��ǧ�7�6���&���A�-C��G��p�(�3�>���ޚ��f�����7�C��S;G�0��:����\�畯���<x=����W��㥇�H�q�N�
�>�Ζi�<�oQc��Y�%���IZ�?`AR4��`w_\D�=���V�v���+�:�âƒm�QE�u�tyx?�z�(��'�0;4��U�;�c{\����'0��{�F��9��?w?�Z�y�ɣ��nMl'P��Ҭ��{��΍�<8Β[HYfs�%�a	&����*����{��YPX���S�!D�����D�P�thBP��Ȳ�G�I���A��??����YUc�2]�a����n��O7|?�K�*��
G�6hL(�wL����h�d�k���7ʢ�.G\S��	�#��Y�x( �9,p�ER<R�˳�ϱ�ڽc�|�10��R�;6�����xb�p�;G�Y�,�V%�7N@Y_sq(I�4��e��.{v>q��8� c��U����o����Qە�c�����u<�9��&Ԕ��1+WxyI�s˽n���|TΩxz�� ;�9ë�����`��]��� ��l�����UuJ��aVA%�m`��FM�q
YѿL��\������x���5"�d��V�Q���Yd|`���F��~*���O4����X�Vl�?W�2��x��U��O;���z�zpf�1E�2[�_�R�����z��i����,% �����D&k�\������j�L��W�`��2^�a��@���v�V�[)^D۬X�$00�SM�I�k��q'�+%C�8�V7�®�'AYn(�D�f�D�p�y1f@�d�C7��K���w�Ϙ��&���d�	/eDR"8$��&+�p��vE-d#�G�I��I����o�H�н�6u���	CS��=̚�	gk��Xz�Zt. ��j9ޅpv@��ôx���%�5��.���$�x�0&�gpr�k_�>����%yt�+���ȽB�{8Q`�sP��+yA�f�~pK���Ϝ�O�V3�-+b�[� ����Qs:�ޡ�ɉ1e���㣬��鴭�����*2nAr^-%v�c��c��2��*�_���n.�A�-�M���IԲYo�1�c�9�f>���8��-��)` BO5dY�Vf ��-��o�D�
m�+J#�|q~ih��+����d!k<���fq�]1r�*�`�#�on������Y�x�Z-�瓕]�$�#o�qrh쨨h��jS�g�6��]e��ΦK�~m�\@y��O�U6'�?�v����@T����<(&��ʤ�̵��JI�����Ɩ��J�:��7�S�n�JD�r��@��{�|5�9��>	� H5]�sv�"���˙�?�kz��]�2�!.J�_@6����������2B'/��t�WN�v��	Os��l9�[��Uf��îK�;��B,v�&�,n��ġ�-qΘT�� �Uځ��	�Aʑ�A����^W��i�y䥇 �4am�(�7X�l���� N2Iǻj���:C`�+��a̸q'<�o�mw�Tg���L�V�<���-i�i�=%+�j�R�C�aۋ�SNWH�~�מ	Q����š���3��Hѷt��;Cۇ����8�����v�
9�3�_�Y@h}]�k�1U	o��BY:-�N_�g����c"��[|A���5qC���q���X#�*�va�{���Om��A�?7��H�����Q���Qf1��|u��Վbs���(�g'm�Z�au�L��V���+��j�쭞&ʎ 뎓�t��kP纼&8aPzf�B�\5����@M�``�9�<��w���.k�{�4Щ����ޏ�8�@9�Ei�1?�z� ~DM}�B:P$̃�"�ɐ%8�t���L��]1�!������L���i��d[��Ǒ>�F-�F�Rz���/{'0�O���a������_�5_(F-a�+0��R)Qܱ+� ��3%g �P��d����,#K�9�Lx�
r&fm�q���bh���u����&���^�*kM<�\49)�5I+S6���@�8�.n+����#P��H.^�a?�Z�$W�B'w$�_'��Y*�Ґ�'����w݀C�ϧ�B�}0��㜠��v�/΄�ͤ@�u��>'���7뭿�k��3�1�D& ��0/���[{B3��۰f"������I-���}~�9��!��������Fl�\첌ڞ�P�5ِ�-��D�q�T\6$���!]v���_e@����E�0��T0���9C�!S �sѥ	�.Yԁ8�~9��"D+�Ukd�5�$�؆sxH�,#T�
y��{B+�/���E�`ݨ�!�mrY��[ ���g4!�c3��^'V>�}T����l�W�9m�}���	�QL�x���/���f�ѻ�Ka����z86)��eA�� �\BW��fb��1����^���k����?�_}����~(�٧����
�r�8r�!F�_��5���oA-�C�HY�n�����\��w.��=���k����^=���CDF�D�����:����OD�*ܼC�M-&,�4�5.җ�u-��-��mg*�����a����U��������5���!R� 
c�ڮ\�	��et�#Ǐ�����'��2�G������b�^Y��&2��[喀K:��Μ��z�|N��?�TH�O�������3�B!�$�#|�7��*��OF#6~����ym0	����Ϥ�.F�IO.Va���Vn�r����:���eX�ٟ�^k	�3At�f��FN�m�iޣ \�yP魑�����S�#0��2k��x��L���zz��~�|e��^�\_"a�U�\4�(_��͙����E��k�V�s�!��D�!3��C��A~?/1�3h��a���SI�v�
��P>�0CĽq����q�K�0�{[�����֘yw1C�^|�\(	����Rx�ƙ6G��� �ӯ[��0h� v��W�y�#�rf��.E��ͪ���b�O�;ۛ+c;vC$k<Of����Q��齥�
((n�z%,��~�LvI���-�a��E<^�N�Z�ek�����F��gI=�~�*�a��A�g�v�������GW��H������|�5�Z�kM�v����)����A	�nb���B�'��S�'��B%�2��`�Kc��6���=̖E��n��k�t���ۻ�Ϡ3�50����q��Y9��~�0��l��1��䆤)��-�(�C�
}H���IGh��0;�`[tEG��=Q�.��X��k/�-6��O��IN��KsD@��a��V�r��@}D|�D;x@ö�d6�)q����=E^�w�L�|�?�tL�e�>�*�&�G��W-=���k��O��E1�ᷕ�ÿ������>���M����IH���҂oz��}�����3҃��9$e�l)��(�1x����(m]]eDde�D�3n;4�͂`��WO.�M�a��-�l���{[���9*��?���7�N>�?8[���������.p���9��3'�5�1�^�0��1�8�U��P�+VAg>p��u$���
�1t�68��*R���>.���@Jߙ�|]~.�CfK5�]�1H�0�����pszB~J`�ma�lgĕ׿{�M��j����_�=[�=N^|WJ�܍v����~dp,	�|��c�ћ�'��	6K)Z�%�xDe��EO�,C�ǆ�PeJL��/��mE"�&�Q�\WqdI'i������ y�ك�L��(T؄��gle�	Al�0��M��l�zwA+�p˦�JM�nN��.&�5'2��ar�>��s�j�������b�֑���i�0���jϻ��pc��O
�3�ۣ/6ۦ���[��}Htj7��e�� }��F��)��3M�ŀ�C7�	֏ɰ`Եʫ�	�.�Z�ۖ�U��TS����VXqDsoa�7E��@��w`SO�7��H��
�!]K�W�� ���L�x�t���!�xY����^!ؖBUtL��[An�)ˤ_<a��t*k����>��;��"��H��_t�j����U���ȺU���+LH��4g�;��@��ǅ�������]��D�(<� /2�Y4��#|���o��B0�(����%�Ɂ��^��tT-z�Ԯ��,� AF�X���-@j��m�rd(�H}�]`�n��(ӏ�%4�m�:O0�	�ݐq�
XM;e��d�P~)M�������OC�Pǡ�:}�6��C��hHf��
�2hn�E2=,����h��t�Ii���#���FTaG�uh�WPi_���(��b��B4S��n��Gg�^!E; �9ǣ0�]�����E?�AB���6��?aA)X����d�.	��"ي s�e��.�����L��x}!�u�CFH0&2�p�<B���{\9@'.A4l=f��8�TxyC<r�M[_���s� �P��9x{�[=~��%�n��đ�>mR~!�J5�V��˦`�|:��/��b�8�rws:���T���M¸�+݈�V�g��ȵ1��^�g�*��gVԱ�n`���E�Q�o+qp"eԲNu���Яf��*�'��[�H׍@V'062�/"$���Uv͈(��q,��̡´�����X��Ja��-�<:I�B7u��KCWКx������:	�b���v�}��+�I
:8����Bυ������Ļb÷������_ei<��Am3Ȉ�xź���p��<�f.���> ($�"j*Hr=�褢��Š��v������ϯ��X�m�x$�i��#�����+OE�p���zX��q$#�j�����zd��Q]E�T�_�eЂR=��5��W*�vz���C�Y��9��q��䌯�R�����tο4��ۋ����d�//������T$W���{ʋ� ���Xp8�)���/9�0yoh��;H�L1�fbuj=s[�*_�s2�q��N�[��>F(s��a�.wĒ�n���}�"��g�ÿ�S7�v�	�����r��"�w}'-oy���*4C�����E�]��H������*�cK�{hy
�5�T@q�.	T�Sc�S��1����)u�ը�ޟ��V��C�e*6�7���Wyܖ���8��l8QՕ�v'��`j��р��XĢ�Dʦzf�u��n'�E�|���/��XRg�m�&Rj����1?sAؙ�f�ON"g�}*3 �0,�z���%��C%;��ӷe�}1���[r�V$OSl��a5�E%�����gW�o�C�`���vc ��.F��t��cBzGN����@V�s�4PO��6�0��e�Jf��N���b���h�:��b�a�F�I����4i����M�>T�I��z�t�j��Z�����N�^�+�.n�Uu!j?T�����% m�6G���#o'����0x��]Nu�
	���t{!qS=W'���u@�$����"��vڸ%��9�2�Z�$|^��*f�jN��NؿF�G�O� ��I�����fp˘�Ԯ�Y��/]�%χ�����eS��G0�{67�ѕ�d�mqc�i�w?�}�ʿ�t'_��( ��[W~Y���ɵt"P�&H�p��O
_iq#�l���.3tIY�+��sAٗ�W�jՉi:J4���S�1_�"!�fF���|�U*;y�Ek:~�<�Zui����<���̘F����a����>�削��d6�#��끛zKɬ�6��W=��25!�����6L9�*�HMG�?���&b	�FI���S�T^��7q*$UV��@7��Տ	�?�E��MQ�N��}��V�l��9y$_�G�c]�.��hP���"B�v�Y=@�a���!�T��I�p���ևXR�'�ƍDK�}���sSE=i,bBo��lֳ�59�S�`��uw��y�ݦl�[�@ޝ�R��D]��6z�f��gSxC� Z$-X����Iq���� Hٳ���Bp+��(}s�)�CQ3O� A���A�2;%��O��o
�X�$vU�4�ݡ�$�P�7V�W���RR��WYjC9ട}'V�+�=��L��
l��C������+�yi^��^%{����!׎�n�3��ʯ0�zKr�ժ���;���R���۽���D}{*�U��Kk���b��`6rR���;��h���Px��f��6fe��$I��	{�}��͢��M�a�#@�yHLҌ��]�*26�v�Q�(����.F%Sg�Ic^!]4�E��_��JH��rm�s���+��,^[�غ6]Kpa%&9�2��������7�n�EzAU��IX�Oa�I1I{�w~��i,��z�8 �ߕ�$�Be]
�f~-�bh'XhR�0R���z��bĹO��!���Sܜ��_ra��6H�; (Y*٤��+��I��t˝�'�E��B�Æ�l�s������n>8Z�3=�D��dJ�K􅞛�S��t�bwX�^wy���ʄ�j�N7�r��{^�]}�0`�5��cn�]9a�z�~7�ǭ�pͯb,-/�l��`�$2͎�纽#:Ŗ��������-{��;S�D�Fi���%�����E��V�j�ӷ�G%�={�����^����J�eR��*�XW��t�]�\Q�ǖ�Y Q*�GD
��{TE��(n�zW�IUZ����;�l����*5r�oʘ�^}	���wlv�"i��N(�)�'�6������Qohy]n*�n�����\�����H��Q`�Ѻ��k�`��	�N��kH���O��v7�0P�C}������J��V�f����s<�s��{+��<�yG�`>Q� ֑k�!�oa���?A߳�`Z*"蠀=yS�* ]X٥���gy4��U*�N	�<5���8�/T4�7�ض@�|�/ϯ`/w)	}F��#n��,{���u�e��1���f���d�lP{g�$�g,��0�_�� }�CD�G!#&�.�/�RV5P8ZL���[�!56�B��Lü\J�Z�`��+"4�B7?�;��qR�w MN�će#胨v}ri�1ӏz�fDw�r�D�U��s�mY�ckTfYZ�HlS��?���f��g' ZAu���@�Ll��qB#m��G�C��_�����}(F௼���q4 ��[U�_DzC�\�D6E�k���Gh�(1Fzx����0�V��ζf$ZN��P=;�`�Eѵj:���=�Z����k:�Js�R��.TTDXm�����^�Z���6`h�L�k����]]�ᚋo���~O�6���1l��6tN;4W���� =�"RhAoʫ}��9�S���Eq�A��
�h}X�����d�&H~-~��Ծ�K��t<z�yI�����n�����\43�'
a>
����W��VKr�r���4�z~�Q��1̩���dP�wT]�w�&,2&��c��6岟|��{H�����CM����̠e�����2�H�b�A�8���+���j�$�vt�_!��S[dF���F;��2,�=�	Ǝ�p=!|gm��+Aa+?_m�/����`Whg�9�f9�)�XC�����JQ����չ-k���G�1�������>�B�|��8vL�C�a�ټAF7*��s
�L�%z�	�4E��kz�z�*��u�U�ӔBb���%��
h����v�P X��~ 
A��g�y��+���8k�*�y�a�O:���f�n^�@Wn�h}mV ��LK��!񊨬\�G͛�M��R𞣭]���CH~y���,���V�e�8}�1��������.��-�?�F��f�\��'�()�H
מ:.š�X� �9U8*x�	���"����^2�&��O�(묒��� ^���N�z�O֬�x���d0�iLqx��$�=d�� ����k�S�V����m��]	$�ފ�!���O�	�[����B}�^s<��j�skV�7�B~�X�ņ��Tp9MKkݘ����'��m�E�t�`W3�q`��y ��MǄ�<a�*���d����r3�n�s�ߤC}҂:���������R%��w�s�-B��<��%�B�sd��������	nu�S�@��.Ms�C��-���?9�\0,��O��U�,_�ɠ��ӑF���\�f���$WE�<�F����i�m8�ǁ�U
�2h�E��Y�3�Yt�IEUD���C}�x�`��H+��bA	���Ŀ&�GB�j��Vkf��V�M,<�.�i�r�`օ|i�j�'�_�����o��V��ˢ!�^�ɝ�J+���\x`Q���A�];�+8�_�>Qfh�:�ľ����2.�1���d|_X��O'j&�>�r�,�n,M���h��'f��6ј��[AXf�q�u2�y�nN�~�eG�Y#Ǿ�A�D���i�=���aD���<���B��u_�V��u�դI�I��(*���Uu��7��NW K�$Ro��J�s��/��ޜ�;P�l��Ժ���j�;���dr��[1���s�+�b}��oG�wp�L"[�v�'c� 7�P⨧�7�q����!��
^@=�!����R�,�
�L4��w�Y+�+�3o�@�&�^0��Ć���o��N� �V�&	_���x�g�a�.9�1!E�x9I�� �ѣ��`*��D.(��8�.��8�	�`2=�b������@@�4Ö��aē��}�QU���g��[|���%VNRW�<�o����$W����<A���)�P�b�3yO�tr�{3�҄"��\9,\��_��+H���l:��녅;9��f�ƀ�AaG2����k,8��5;7%�,�e��G�?sH`��k+ B���.�z�ۺ{�`���A�� G��B�T�5�c��;���n�)]>��*kjZK��FQ���s�+��h?�u&u���l8خ��ˮ6�ftyח�����en�ҵ+D�	w��n�D5�nkZQ����5-gxh�s�#"vn�����W1x��H�����Q-}�rk��uِ�� 黴����8V��:6������`�v�����/�6N����0bh6�{W�I<��]0��Z->�O?ęL��r
��Oz������\'4	(���Z�ߖ�S��6�]tr+������62F��715�z���_�ڸ�?D����]uh)�B���6�f�(��X��qT�1�n�E�e5�Tփ�r��g��X�{���2�8�s�������T�,>�Ǫ^^镫�X��y���R��8G,��K���5�<f�����7=ʑ}�	�I,��H�RCEph}59T�<yvW�o+�SMS(�\�K�[���C������?&�� 4� ~+�6�7�=�)��|�O%�+���p�d����+�uZT:�Z��1uV;}�(w� ��7:�τ�=�oY��n��^�o��J�����XLTläAO�Dy=���M����E�n��!�����"��fɒ��aIXϏ�[����%����-5��Qxt�_�U���l���$�·�A�4��+�.�I���;oQ������lￎ<���o۟���c:ss�Դ�me5<�����$K@0��Q#��G�w���6��T��C�.�|���F6�;j���g�z�D�|�T�n!�c��_����"۾y��e�.��.tIL�Rt&;��0m�c�m��/I��1���I�wBl�t �6mEV������vO��kՈ�L��Ng�/�\Õ{#��$���&vAeM�L�E� ��=g5y|#�s�xH��y�v͖[�p��Yv�$I��VEom�Q��D��詽���5 ~��C��%�s+)%,�b,"W+j83��5��t���:h��we���46y�D�'{#�����d+͠(j�}>�.-��bp�bz��6ن:N,F^�M�0jL7��[��\��|�G�6�ä�E�d��!�j�V�4˽��cUٴ-�c�_�J��E��8��\��Z�R�b��ls��!�W�/�G)X�=�Nw��])�ݐ]���pΩF��$�u���#�����H�0��0aW���ws p�ާ)m�������Y9�\���Nsza��)u��s����V������-�����ރ�9�-�����nn�9�g.6��gC�'���cq��]/����a�#I&�Y����S�����v�5�<����"�_�u�o�"��
4�s{�04�r �4��

l�%,?�0�^�M����*뱆�M�Xy�E���}r+����̥W��x���F����">iV�����Jۚ:��l��Ȩ��j:�V�_���l�,�z���������s���@��v���Ֆ��o��U8|W�%C���E��u�姮����~�4lʍ�D$9 ���D�i�!�>k�أ���r�g �Ñ�Qoi.��G�8��s�Q�i��JWi4[PB�X2�ǴE�A+�d����:#<���Y�+g�&�7%�(�U2+�\
=�k�=S��}I�w B�R�L'���&������wp1./.\z���#w�Ӑ�^��KC��9֗6���A|��iJA9�� �k<e�)b�]�{?��~O��O2z�����B��(V�j���/d�ZL�{o��Kc�ѰI�n��;�����[w�kC�nc\U}S�-B�/�.  ^[���[ �b�o�C�)�?�*ۅ���.M�TV�l�Rx����zp����Q(��t�]b�:ݐ��R ��hw�7��/č�$[m^�>�D�����M�fu�ɘ�z(
�h��[��6V_5���v��JC�>'0�+��c���� C�U���)9s��i�׼���P�k���@d����*X�r�{��s�=
۫!����C���#;��g�-�X�\����$�@"�7h�pI�)a2y\�L'��2(�����J>h���`y��+������^(a�f���Ll����:���G�C��A�L0�����Y�d����rq�q�|y˻�kk�g�f6�ah�R�vG����?���o@��ʴ�K���v�U�j-���A�s�r�����H��ʻ2ּќ'�dY|�r+Ɵ;�pJ�d���04EW�.���H�.:8K	��7�G�P��f	�;�|t�p=�7�WX��S���`+]?�1WRߩu����+8�QU���pi}^-�8��i�c�F\̞�;�������H<}3�ԄY��8�q��m�{�p���ɒ[a�Ym�3����<��E�n��@8����f�ב��� [��ZH/"0Q�g T�I��:� W��V 7ypp�R���8m��˩KR�}���J��^��R M�f�[�~�� ���t�G��X�BlN��͝�=�L�{��2z�]��u�!��`n������Jۃ(�Z�w/wb��J��o����}mŦL�U�J �GB��ށ��Zw���6�ZY"���������c~��N!�7�=$�&�`̤/�e���S�O�i7�� �χVo?�ыנ�\�:����RU�)��|��9�I�a�X�E�����?ٜ�D��?M8�Ywe��s�"��WgT��N�΄5�W�m��Z$8�@�h�W�D�&U�`��D�oBO/��wJO���و�@����ItT�������;�a}�L����j|�@��wS�O-�����>f��<��.����"{�%�@�����/m�7:�6_�c:!RF|w�/0�h:��ZE�0�2��ρ�*v]�H�����n@�	�?H��?CP�hԁ9J$F������I�9�D,�i|8A��^�>>"lʇ����e�]�X -��@�����7�.b�}�^�_j���O[�q�DKR�=LbY�!��j��!�XT���/��;H���^@|�lv�����%���X�
�ѧk��QQ�̼����f�B]d�J�sR��_�ӽ ��zS�~p��X�e�k�j&󄿨qO��y��S�+�A'ss4���*Svc(���\���Lxd�^�ӣ4`�0im �I��0�׳w����x>�e���ȋ#~^�N�����F{�2*�P1��1|&��F�%/T��J#�m�B'�X}�z��ޫ�B1���q���h���	�VC"�	���U~cq�2��ոd\�EIn;���ծ'�S�l��G�G@���n�@�N[7$:8���K~��B���Tyv��V���V���r�M%�5�`� P���Ph�P����w�	�Ľ�֟��O�l�ӧ�{@�"��^pB암��Y������Bz���k F]q"����g���gb�;�L= ��:���'}3�J`\1�U]
�j�2���c�%��S�ώ�>2vKj�`�gte������u��� P)UU_`�Qr��JZ�r�{�tw�z��	|��h�G�f� @� ϶�6�:\��ݫ�/�WXd�3��el�E��u���kr2M�����k�z���5L!��(���SbEcn�'�ۼ���Wy�=��/�^|��O6�X�����a���_Y�!Sk��F3G��4�����0k�́Fޝ a���:g���.6��2��{�N�#�3?�.~�h�,s��p�u!N��H�P�:��-�)�t1�9D�+s�)$7�!�5oԡ�E>^���W&o�D�`��%ҧ��7�D��IC��]s�	�0.{�h	����9�i�Q���Э=Q�u��OA��(!GA��V��4`��JXz�K6$��%���j�Y������J�Hۥ�p���]�0r���y>f����o� �m	�n��k�ܯ]<�V�x9�Kv��< ��MWU�+ܬ������l�-�G��NQ��v�3⎺eɆN�S���>�����@�r$G�%<^�ur:��*�zu*���� ۶]�u������69�J�b�q��v�5&��1d�����{|�� ����9��H>���H�|8���!1m�̖�KI!R�ނ^0�&�Y)�����5v�zD��)J�m$��Uu��C&��!y�f��z�?�(@d1x��/�w$�)����Ej���͇�K*�/����F֜6i*���w�KG�)�s0-P[�N5�&vF��޵�5���5�/�Rí�fKz�5j���˩�U=`Gg[{;����X�k�eep�`�2�7`ph��������xA���}�P���W���4��<��l<���qy�+)��z�?Eo���R�7[ui��_�D-��1� ��{^i�:���Yj��\_�-d��F5���Ę��O�Þݜn�HH���AH&�MT�	����ۗ��[��֕���U� �W+�L�s�(?�g�N�Gl����5-P�ݶ�ۇY��K'ᖓ��YD���F���'��.���-�"{�@=�rėFo�/�[��t�m6�Q��`��!�����Uo�Lb�S��������A��T���䨕�������t�u��d`����t���J ���e�>���¼A�� �9�
P�ԓ��VB����)�[�퀺	2eV��w�${�ܷ�Z�St�:H'�����d(���i�6�J�H�o8{�U�x���Ƒ��< ��i낏�@�9[��m,F��`ȃ��1��P$cZ��%5.��闋�̣��Ƕa�Y����X\ϻ���z�g�F�p=+��K�������i?CFDS.���o�qY:�w��a2v��e&��	����+��ƼJࢅ�`@�X�LXR�i�M!��cqP�wX����L0'�����
�sf$~��~͐�:���b��t��a[�磔4��L�d���=��Y��|To�D�S�v�>d�D|�MLP�eo�M\z�h�V�R|�7�Yp�[2քU�(k>K�b��a�f�=]W���	0Z�JY+�Y-��f���C����%�tS|oU$�+~R*�cvV��F[��#D�N�U4�8�����Ε��thQ�Y[ہ�:v���5�~��#���Q':>ך����<=3����j3�z���m�\�x���S�[�Z�k�w�����s!�?b��k��͙AiK�G�� ��5�_�ݡ��M�0W�S�r=ਦ0M!������9p����N�E���,e��|x��6Gs����Q4����C��HR���_�1?�6���o[�8����x���c��M �[o?[M�2�*Æ̈́|g�uS�����DƹBQ�b��פm��T\��ޕc�����ӋR�`D���IV��^��(����������Ci�w��f�\��[�5��$gB���_Ah���Urk*�8����Tg��d�Z�hI�� ���1�;h����ɢQʤ��6u�Ô65�9�p;wlz��kf��� a�1V���L��(��b�U�,~^�, 
W^斓~��n�k��d��I�u6ݦ��!�")\��pQ ^��=��U�����ve�yB��U�L��V����*$Q��l�qFmYx�\��w���V�j�I?�ƥOEA��g+�+|�J���C$�}��_�C� n.�&�,��`[�!�S���d擒K�s�$̟UO��y�G�9G5�"&\�S]6��>w���d�����[�d�-r<�l	ّZ
ܴ����Hإե5˕���u�Q���{���؎h86�o}��7L�C�����a �(/��
a��7�����2�Z���L�G�]^]�m�$1��N�"sW�\F۪UJf�dT�)aR �6V���W�cԙA_'�|�>c�8�ٝm�,��D^���Ǚ��y_����p��Ca����y
�+�/����m�h3��޻X1��U�A���� ����G��Q�7��@ǲ�Nrh����P��B�z��+���/d��2���W�:�c�����W����48�͕F�`��g���L��Q6�L+�8���],S��1�6�MM���� _�lަc�ԆNR���+���P�p�*��]@�qG:�j�SWGZ�vϬQ�{9$�e���vnAt�l�)�r�Yt1�jHG6�5�R�y&�|9�����%(����9g��]�I����<zӒ��)���Wf �=7�+k�c�.4+�PG*Fb����)ؙ��>��	�\m���}� �S&-��\q��q!<!g��[�z�/d�<Ru.�������J�@e��~��4�]S#�4v,�[}�rBF��>���D�0���`7�!q���S�M�M�Gٟ�&�)+@�*Uw�<���+�7>v���Xt'/m��*7�������< �2|���/���K���GB���4�0E��'x�����vE�����]�������~����@�K9��&k�S+.��1��S��Op:tF�f��u�����@�
r*D���3F��<E��(XG}���W2����4��?gq�!X7�Mjk�0��&�)`"RM��)�c\)��8p�E'g�VԿr�݉*i^ؒ+�5+�TN4��
�D"�E��-ߴ�ggZ�\�u﷑� ��IG#^�ǔ��ai���.�C��pYxuW�!<"t�=���:���ҍ���Ƚ���T���FhU�1�����Ϩ��_@�q�mK]����9��,�^qRٻ�H�YtEz�xs �L���h�_g�� �go��w�m$b��_�[!y��Q��T��T}%���-��(�wuJ_$���$`�Y�K��;��ԏZ �-�ՆT>C�u�
6#Uc���yr.3�l��^��Av�)'����:2�3���v�Ӎ�jlE.c[ :�>�-�����e㯌�jai�l��,Q�/G@��S�/m�QI����n/���a���rD��X�!
�vs�<(��ڬ־�_i_���Z���=QŅK]	��լ��n��l�H�*(,#��5�)ãJ��$��H\�?9�mS�u�J�
��G��5��0W��8�1�{��Y�v��@�*���9��Y��%�_��o��mjHV�X�<6�q�0FMD�,; ����)r��U�4��h�)� p����n��0Ͳ����`��h#�>��Y+x�f��w�$}�����F���|����'
�,,q�('���O@o���ڣ�\�¨�Gn�2/�/nDR�x�xo}k�|%S�"�_{)~�	K~d�k�,�*I4��E��WKY��u���f=�i����,�[��RU��Rm�!�X7�X��������v���qW�l�Ǟ���6�����V�e�։�+v����xl���*p�>��D4��3���z#���@����KL��!ۋAMq,�ט6�W̍!%mO��m�(&U{���70�V��P���{��F�z��/t�lk�W	�B�y�n�����#�}I��)���,dP_�h2�l��rs�bJ�V�T����%�3+��.�|��0�End�

�����~�W@���x騯S�W֘H���@YyiU��:*�a��%Ta�z�q@�Q�p����P��oe�[,iJ���|�7N^��y�Qۨ'���^��p�����$��-��8#_�Ҧ~PA� g�ט�sTѺ�
x�>�L0uY����HA�㞆�v/&���ԑ-	�ℎe�	�570u3�9)Q�|OS	Mp���s�R��Tq�!=�E�P���0\)J��sԏϻ]�v�����~"1�06���%�o�G�ʹy}?�uyQ��_1�q�y�[i�0�Z'[�(V�	�>��T�`bk���޳���[��T����rΏ�<e6o���,���ð�BK����NIz7R�A
u̥V2z
O8rO�2)[���A�?�_��W��(sD𿷢�)�V�{�����+l�q�|��ʬ�-�%�ZN�Ea��zXk��^j!��e�AA���~Z�d����Dw���pk��Fێ�Xh�u:t��*k���,Ј(d�'rfWh@j�",<�t̴�_���x�B,v1���vͮJ�ǐL։��B��6��<g]Z�W�3&e����M�1��$GGgnL�r�A����|n���������`����G8@4�wB�'H�z�<�0��_&�N��a����n>�z&=!�G�/6*��?T���<*�Bx�|�!s�~�[����WG��|�AW��7��!}/��H�B�����X�b���e�Um�v�.Q)�e#u�Q��ѐh��e�8�i��D�4Re7@E$"H+�>�l�ۖ��.���>y��`Z�4�/���'�RT~6�Us������hnc �׆f zV���:xZ���ygB��a��>��(F�Yべ��td�O�Ň,c�F�1"R��rfZ�E�DӠ�#|Z��}5���'C(/��Z� F t,��O2����R�Ȃt��/K䶃�]���8D�!x��f��}���f�}��g5��
��\�Ȝ^�:o�oK߹(����$7����l��� ��H .ݳ���N5����y�C�}D=�;!�7x�'��43���s!��3��⸙�I�ͼ��|�H���yvl�Ь3f�X���۪���@7̖W!�"C`{V��k9�,��o	C[�K�-_��[�%�g�b�͈��D༢��A����
�5i.=��.v�-H�ɆFUi�k+���7����1IK�!�~�}*⇽��R��!����4q ������_�M�n
l���� ��ZF��Ǣ;8���@P��Q0�Y���w��G��Ș$�WRH�����+����r��"��F�s�P���O���P�4���K�U��_a{ձ'z�fzD�9o��6��%��+�����*�S ���X+�jE�a;����R���� ��,jO�Q�<`SM�y�<� ^���sw"�kC��X��ƅ~ȝ���%�O�}��Ǵ�wJ�@��*!����{��e�4c�7H���]�w6 ��ý�(ݍ�CD������OX�hèA�#�n|�G~W8�M3��.\G#q��α���:Z��T��m�H�@��34����;n�uu?-
0H�KI�8���2�f5-�w���n���}�Y�r�K��u�+��5������]�K">ب���J��0X�=��xǢ������}��D!�S��K��ϻظ���q�u��m��E%mJ⸸�R�y$�� g̰:��]ľb/o����6�7�^��Ouok����������kz0q�g�`�Փ׻�P�F>�����.��F�O-hw���4��s
��>����$�o���.mO]J-G�s�E��(���^H��cg��J�<G�|o���~��I�n�Mﻕ���D�a��M��j�����w�n	�	����:�_�f^��)�(�P��e�n�{�7�JE5>(`Z��g:\�6��5G���TUC�P�C�S�&�Yg���#9\�{t�"�\�N~`j	�J�h�;��#G���"�q�D�&/���܏	J.�����ʤa�;�y!���w�k�"M�2�SKt�)�В������9^!�J٢o�%��e�	 Z�jISѯzÔ������@�=�)�:� 5T�`�f��HRU�@������ }�`Ë_Q��n.=`~���L��$��,w�!�jqt/>��^�tr:�[k]Q��+��+��qt1���H���W�u.`��F]��
t#K����}���T����;��g�E�5��w��G���8�4�1h��O]ڂ��{H�~S���.�HG%1
��B/��{%�H�J��Ǖ��z}_p�����*�N��GV	r!�v��q�r@�eu��I���1��{���`��Q������|�[�Eq�L�e�w�U�̺0���rg��祾@dCK2!b"���]���ч��6�g<DE���d�����4�o�kq��;5J΄��5�]B�ģD�P�t%ސ��!@�s�����J��_P\ϻ�QF��g��"�n���ˮN3p�On��5��MY_�3�M|�i])��
(Rh�h����7�X7�����v"p�!���[y��N�Q��덖Gm�!%�t��/aM���y���i@�͚߫F@��!0��y��S:LKSHlX���f�/��-��n#)bYU�����H���3!�&w*$P&�\�3Zi���$o��_��;t��`.M�  ��y�WrȄY`��jdЯx�s����rY�V��
3��KKċ��9��26�_&���o�.�^��S[ՠg�w���R��l**�ViKjb��ǘ��`䄸��� ��:�E$�#b�\Q$� g��SEWN�ʫ��$����MMI�6 ?�y���D��"�R�tX�� �f�b�j���������T���"��2��(|���`���z���G9.i[�6cqC���V��aKl�)�^X�*�G�8��7��׻;#����/�P�?�4�EV$q������TV�(Q�V��ӈ����Ī��ч�Ͻ�ȡ�r�Lh������~�6�Ñf!�t�[u���-�}�+���O�E��#�(���k
:P�`a&hտ�#�g8��W�B����j�}���ϣXJ�����5�dL8�耧�:����,���#�~\�o��{R��*��}�H8�ʁ.��Jju�T�n�j�a�*�oc%�Ċ��I�?��lA:�4a��u����+��1���XO:o$�{�
�c���Iܨ�j&��xY��/Կ�׫5�x���ܛ�鱣[>l��cN��=���4b���9�ļ����U$5��1��d�_�^�����=i�
��pF������C�iiL�µE@��+V۱���8�bdG�T�i� ��{�i���%��.T����ws9��H���+@TTx'�����w��\e*$�qB������g�U��g��Ǝ�,��ߕ����A���S*�ٞ��
�����9yj/i/�tt=3远;z1#G�<[(�Gy��2 ����z�W�DH*�oR�J�>���2b�b8�
7IOXC,�J�6��3j�~j��.�x�c�^zfc��J=�5�	�`<�uڟ�_���Զ���탪��w��e.�T�Q���ZΈx <(��� &ˌ���R?�^����O���ѳ#�����V�mZ��ϭ&H�U\?O>�v�H�>�j9k��+�6��u� ������U_��K�tl?˔uAs�g)����z��q<��o#$'YG���.�u��/��fw�~�kA6��˒m�y��2��h��ٍ1��`�K:��[�AO`�B�I�ǖՆ&�G#��?�������J�r��y��mn��nj���V���7f�(��5V^����^�V��/�3���z>�!@Zy��r��Ʃơ4��t �:�2}/�9A�QH���a���>���,�n*7e�7)���C��6qh��a۸��?�`|���BX�7$�6�=�\�(ë���j=��GK$e�9p�H�R�z�G��IDR>7��K޺I����m��(�u�,g����t�������;�C�w���ρ�L���ż��k_Q�҉oa�h���&�G��W�O�5�	�n�G�ޒo�äO���h���G8��n�6d����ȶ6,��$AJv(�d4�N�j���u��\����7$���0����)�@ >atHw�&K]N��D�\	��� ��(����̽k4䥨R�,�wO���\ ��5-���OW@�c�����u�R�&7w�#��$�N!��=r�U[fX�Ln!�4��g!9\��J��EZ�����asl 7A0Z���wP��zl4���De8Rldz���>* W�P8> ���|����>aaj�T��ʛ �B);��w��w����$���u���_����w�,!���Q�ֆW 7*/�Ka��F�Z�PL�%P>�%���x�����h��x��?fz��ϻ�>3/v]_w�o5��AF�R#������+�ZA��x���	��f��e>?'���C��V��7�+��T
��#8=@�P�|�O�սJ\	��7�/�����*tA�>s�$q�wXt��4����/�	}�UPO��r/����t�(TG���rK�@�[B����;�ڤ���l���A7�='��&Y���;m����+fR��<��v�9��掴x1��n�&�6����H�M(|羽t��5�n��RL�7���==ЮM�5OXQYDkn/31�)N���i�h5��C��2�����"�r���I�O�R�h֛Qi�P��'	����BϧQD�C�qm�%ǔ'oXCܒ�͇���D�\��v�Lʩ��浉~4��U7�>�YJs��؄�6'��2+�9�ƛ���k�����^?��7��<J?l& m�!R��$?�L�cq��B��[���^��hV҃t+7EA��I{���T�/���h�W.���c��\ҽz�i��:�c��*�
@�?��*�j����g��׾��	��w�"L�Q8AzMT�Y��� rT�l�;��*�~w8�������S�e,�h�-֤�e�w)7����dg�%ïL��!ĭ\����	������A�@
���t�gQ��,*Rhud�V������������΃v�&�#��t�M��s����>�@�la�ԐG.#��x��:�պ;���鰏#X;'����<�PQ�+��L¨SMټ���F�a��1���n6�	�8�[4��~���n���ܯ�-нX����mv��I�*%s�Q'"�#c��d�	91��^�b����U=q��4K�(��"gj��=�@c`^v"���{^�X/f��B�Ѐ���m�;�C9Z�Qj��q4p���H>�Cֆ�P~	�:�n�e�y#�<�,\�E�|֨Q���EDI�2qnP%۾�qN9+#�a�T�P���� �	l�k{:F�v
�1���(
���9���ns��$���O�)���.l_J��X��V�.���2�VU$�Qj;���~��$�e���m�g��Ŗ��sY!4=W�w�^��7ǋg+�}��UT�' �x�?$��.��vކ���nG���9�c���.�	q!��/�E�s@��&���+�0ף�iua tG����9 ��C��?`�`�Zw�ߨ��VX��$G5�1i�N��9�+�&�2)HY�D����Ρ�����(E�kL�hU�̹�s]���z�X$��q���k��磕�!�y���;��s�����-gN\*O�
xO)݅X�N!	�m��(<�Cњ�Փ5B���)��Tn�붐�LV���q�Э�4?q��3d�� v�(��m�B���^�R��rh�?��͏'c