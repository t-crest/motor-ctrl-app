��/  �x�Iay�g��\]�9�۹��X��Px;��7�D_���z-{����gN��2�G�E �v�TO��Y>�Sip����ZZFC`�π��	Q�X��ӳR`��sj%'R��G%�yv/�Ҧ����������w_��@w�Q3^�%b|)�A��$�^��<�J���6�����֕��**�4�`74$�xe�#]k�<DT�=�� �M�-ΓS�=��w�ėo��7���7����r�2_o�DN��E�����,
�2m�hSG�N�k�
�c�v���s�5T�[�TrL��(ֆ��%�Q��M��=��,�T�	��)�\���H�`қ!�b�cs׊��r,��QJeUy����+~�b0i9]��d��CÂ�v�����`8L�2:-_�#�@Ǌ�6�I����`C���)�"l�%
�|�պ��}�&�Q�n���s~��#���iC�ulPX�k9Ȅ����0e���^o��WE����;K�Xu�wBZ�pny���nz�.��߄)�Vg�
�UJP��}�0�Y4�Cr�qt0e�.�5�<́y���*�D��Y ϋ	Q?9'z��Z��`�4�95v��n�ܻ��N�%�����)�fL�W��'���^}N��a�D���H�W�g*���2J�^8׻�<-\/��n��T�{�9sAB�&��x�$��A��8[����j���c��i��#y���]v�k�Q"��Y���s�u�ͥ־$>w&�Ҧ��mZ�����:�R8���?���"�guf����WC�+��z��j�W��F0��5!�G����oO���7�b��k��n�L����xdv�W�
���yx����p_ͭ0�*dTm䄾���!�B>9�y_j�v_p�-O�=#2u��v@R�W:\(�z��#��j(����[ �9�*����!�w;MCN�b�s5��j+}�?��|L\���	�B �e��[j`&��yTN��/�{�����Ȥ��	�v�܌�)݉9S�x?�� �8NI�˯B �bTۚ5��i�h�.���3L5�Z���*Ag��%%�<���EN~D��ʖx4�2-��ՇZ�Hӯ�DGg����?��}�̔�R�~�۵t���%��sEͬ!J����ﭮ�M�Tm�r�uw蓠���=���K9RP��'�|� ���-�[�qI_�N�LC_�L�R)�G[K���a?HNT�/����m^�32m����_�c�^�%�� �y���䬾���ո��i��dK�`�6Y(��W"?gG���T�`�$�rMP&��y��9�ɯ��ԧ8h�ZC56��!Y�À�@�xjl���A�����DWco���V�ռ����g'�E��Fq�[�FD��U�҇S�/'S}�y�{�~�!������9Q��{�b��n6�J�� w���v%ڎ%*Sxa�g���D�_�Á�0�� K�C �m:��|��@A
4� (�2Jj_��j#�$M��eЫr�a^K�x���Y�����^�K`��5j���$�BZ��.��؛d�N/����]�x�o@�7��!��e��tt����w{�.���BŃ���;�6�O����"9-�
�[t�F��������mT$�)c���:'�_���!�M�@>������O�J*���N$*�Kt�ĤVc��,�-�]�$��j��d������'�[nR#�En6����n�+�T���V�CŊl
4