��/  ȜNq{�'��˔���9[V�D*��u�A�:t��e�.���v�
*�@��B�x�O�:.� ]�g���1��s�7��}Sb�h%�g��y���)|;Y0r"�z�}�d�*�0^8���;l^\L������!M����.���/�Q?�� �Ob��K>�����۞e��P-@������S��B�F����i�J��I.'�;��2����/9�0��@U��c�bI�����@�!�7�{�[��z���N�
�>�����8G��º�	�,��������@�q� r�*�!�7�+!�8���t<S�j����[C����~;!e�s�Lm�{�Q�h�/S��~�Ԣ^�J^�e��xC'r�&�؂،�Y����gTɄ"d��Ӑ�#r*�߮aMF����z��E'��T��PzG�o�!*+�ȫ|V�,+�#�q�G��~B�.����/깻�!/Q��F}#o�F�����Ζ@D�*K�N��CO]�4J��69�Zr�G;7y;(��ǋ�o4�}|�K�iW�1���������J ��T17�g������G81�~|+HD |�z�x�/>٧B�$Dc�qh�o�C�O,�0��JÄ�~��	���b�8ښ���ԇS��A�9��x�ආ3�a.2FE��;2�#6���
��0j�K�$�?��8֒J����6���p��:8}�0��m��!�p� R*rL�
`�M�9E	���j\�Y�b����K���m���	�����JRWN4H:�%�&�| �������>�c�:C�_!��H��sF��%�JUԕ�,y��3��o��㚆k��+��f"�!Y����8n���b���i:}�����y]?M�W:�/��r`�g�oZ�������f	��'��)�|�S����HT�����ӓc��瘍[��Y���e�%�W;��9�;��n 9{� �h>[=2G�e���%����'��?� ��jc6�^����Vca�
Z=��Ƚ��auY�%���>s�(`�)F5ǒ��(�hl�+F.�jV��ߧ��	��V`=>��
�|Ѽ��J�5־T�FYe���]jGӔ&�!uk{K�'�XoyvxIl�
̴�3���f@�Y������k7htmX�� �m�������Q����Xq�C48ԏx�-řg�B��������e���	�,٪(�bǟ(a1��/��,`z�|�vJn/3K�D�t6�cZ�Lc���`��<����]��X�pEDKƤ������#�~�|���{:��C�)�ht�ת� 03�6S�.��I���A�\�w�$�O0-"-T�q2��ɪU�Iv\�O��ŕ�c�WVY�ΑzR���4�Q�XR?���w�c� w�L{W1؟'�Y޼	��>\(���V�j����g?���o~:����
Q�N�4=%��=K�z�h�����6�6����I�]�]~���`��%{8�s��sO�L�º1e�VpB��ˠ!�u\BʬK�wU�T���FGt�u��cT�2�F�v��b�:�*�!ce-��*�S��>�D�?7z��8Ɏ\C>��_z���"�b:ղ%�sVg�;<�ѵUV�Ρؗ;�`����b�+Y��d�ʵ�%�5�@��^_����ӽ,׹��]*�[%�n�S����݃�9W�W�� �A��(�h�P�w�u-w��7�j�����v��]�t,c���v�N߮���x�98���J�&���56��w�Ԁ=�Zu��Xv�O�l
�Ԉ�,�N�u���QY@�}��@u����qE�)zK'A���Z|%����m���rDK�?g �3��~
㩠�ȋ�ѓ�k\��;���"0uj��b<<ٹ��;�3B��i�d�3��Z��T��\�H���9Y�ۃ�?V�I���т��x�^1���J�S�] #r8�Q�>B`�`���ii�d91	��?�~����0�*ͥ�Gf� ��~-b�'�Ö�`��܇u*Vx�;��عH��O4�h��d`��̋߻GK�����L��i/�(�S=衻�GA���F������.o-1�ܶ1��{��rF?����5�g^�1a.,�����Q�tK��Ę�s��N9���t�aY�!0%zj�y��<�Q�F��W܎Ҕα�~�����A��=���@~�_�
f�>�cV"�u�3f��J�|͒c�N�s"�Z�L0�̎���:a;��@�_�^�p��y:�7� 2/�\O�Y��:�b2ۑh�"Z�������|9���p��x_�H�C�1z-ֲM�s�0�둬,�͚c�TLW������+j��'�  Wg���ڜ����UE:C(�%bf�F'��:���@%�s�aq|=������&�@S�-e����m0�Wf�����3^j�\^~�v�I���m�
�w�~��
	��j�?�"������E���O	m�yF����)$& DHi`V��~O�K0�7kݷ	�e�������V��խ���ʖ4�}���t��h��\C����(��ؐm�:�--�6I��^�q5ʝzu�1!�A�M�`�2�����4y�zE�}C.k`�J�%;�y����[�������Am'V�:6�R�
f��vZ�e�j(���
��!o�?czah�죎�!��,M�o6�$�=���tpy�Z-�EY�*��(�F_�i'S8[����Tys�/��,�/!2q�Ïk�86z�.��"{�͉��w-�P7X�^ֺI&\n�A�r����<�}bZC\}���U��	1[�Q��%Xj�2�=~���T��	�=�� |m�؅��}����@:����}m�"��fs�==a�2}6(�+��##�~y6s��i~�'�GZq�����,�A�Fl�BW�
#�:���1ٷinc��nՍ��d!�!����-ֽ�ȉ��7�x�%�_�w�� Jj3�/W��Y19,��L��!P-^CѢYE-P{��)3��%3��az�ݿ�`�3��(�m�"�ˬ	9�H��5UX��v�.�D����uU�-k�#ssi�x�����֢������=,{�w�:|QC���!�nt�eFIF���_X^�J[p|
X�Ңc=�}ϫ���������|lv5 ��[���iF��	��X��oXgu<�;ŧ	���ml(M�����%�v9�m��_{� 2f�f��	��-o.�E���.ZEwkg�{E*�P�Ǝ���*��������C\���7ׁ�g�>�������a::0�ҏ/��0�p���zh�a@m�՘�8<x��E��s�VdK �����������O�wB1���-W��`�w���[I��5�In`���b��P�t��WK��� &�A6�@��]�t��OXU�Ҙ�s��ApOg�3��zbc�\�ٜg̊`���|vk�㛑�K��ځ֖��!'��?�&Y��0���蚽7l�9N2q�����Bw�-��c��㭉�¡J6�4�̥�fNߑE�_��Dw��ٛN��T�UN] 6��qR����PU�?�xc����詫�Wp�h��ԁP���Fx�]��8����x��f��x���,ꥨ]��&0t�9�Z,�ъ9�@���ҹE�E�6�s�L�����$e�=���x>�\��+%S����mʢ�V��]ޯm�����R�Fs�U��T��i��::&�q>,�Me���:�
m��0�V�� ����)Y�65#	�N<�����W]�2���Ko~ \��?���G�~��fN�rUs\��Vde�>C$�'�Zhc��Ԑ��\�H(U�*o~�!0���0�]A�S�vpfؤ=̕2M|ZC��X���?u�J�� �w��ƚ1Ls�|(�)��v�fZ�\���S�iE�F�ک��'��-��
��Oh>��`�>�*��$���.��h�N��;G��Ǧ+�(�E����ѕ�to21kP�Ez/`^�^R�E���T�SU�v��Cϸ 7�v���;y�3y�]�Wn�YkwֶQ��aWU���!t�兝��O,d�������"��	]���-�=�I3�6'*ץ�g�����\PBaZ9��!@pr
�JV{������F|'L��cu8�c�RI��྄3(f ߣ���U#�[��������� 3ȎQה*��[HA��G���|v>�YeIq)�+�*+�U]�͏U���{V���4���Wb��B_P�ɤm��ď:kf2aI���]��O�f^@$ZV^;��i������)��+��@�T��qA51�:;�x�lG���M����M�C[@D�C�QoP�%Uy�m?X�xv�7�	s�CO^����o��f�]<�l#�Bh��R�����ވ�0��~ce���_i1�0��yB�×�a◅��,V���,3zO�����4x֏#�d[[Ȉ��	���������Hf��r�1^����l|/XfY+�&�lw���\������\������L��O�a�@�]��D b��NVx�� �Z��V#'��5�ŉ�9 zq�җ��@��״�������x��V�m}C �<ż=/�m��b]��ƾ`f2C���F�$1{2t���zz�{6�� {�ց������uE�m���T����.�nVJ�.�?�����w&�O7��]��oI�/�8��y=�VLjg$45C�D(�wm����'���S���<��s��]�	ӐE��L�Y����RũJ�����̯�F�/��-�`v|�4b��<XJq���a��bYQB�&N%du�ѯ��Zsr���s0L�a�a�t���\X-�n'ƺ�Y9oYt��5�?Fy�	K�/�%A�>H�J�A>!9n�����gv�p]�-pr�39��L	��T1���G�Xk�ύD�����2�E���2\N��uFm* �<!̸���u&��b��o����B�u5o`'�FoPO�ΐ&u5"E8���7ir0�ټ�Z��/�dju�>R�&�>j\�*��Q��(X.<>5W��8<n/fU��1M%�%��L��#��=�) ������
���Tw_�V (=�duK$� ��-�(J}�c���?�ҧU��Gi��.�.o�����,x g�ȝ4�m�0M�[7]=R�Ű��
��H�	:Oz����b&b/�?�F��F��Y��o��e�����;�L3����
�T_nN^֬Km�7K3�'����{7	gv^�WG�	$�o^>Я�"���1l�BS���Yx܍%���;N" �kT������c
�Dx�D	�R@�vV�ݗIn}ɶ��֛��8���mi_�_ V�&B�oB�Y��R��p<l��F��jl��ٹ��6H(�^�u;b��s��?�[�2U�*�z�5�U'��e������_��s�]��U�d��!��V7}�ܴjJ$M�7�β���h�qev;l6�&��@˂|�&��e^c�q��SR
F!��]��u}v��L������¥L6S�����P� 6�(�4� �����'�r�ձ��2��M�[�lO^�������3���[*ѓ��;�q��*�-g�Hj$*|����8v�%:��4���6�"r~��0�kz��������<�<ۥdx �tP1��2%��{�g�.;[G�R�3l�
s�d������aׂi��tg�C�8�N<������q�`^n��+��(u�#�Y���p���˖�,�.�G��5��9�0���Q^��c^p� �a5��,x���.�ϭ)@��8?J��?��W1�Gg.���"{��ȶt�ǣz�*Nx��7�����X?�ElkbD�3;^ن�gD���t�`cؔ�� S�z��#��6.��G��w�V�-f_��~�]�� ���U�r��݁L'Z�u�/�_�Ʌ�p����F�_��JLs��zT0b�S
h�5=���LD���~s�Ć�g�I��;�rK�Q������<�:Į���^���oZ J1�X�\ve�;��+�]��f��f&#��nՏ�;��}�׎���߳�'��9�,Q�E�R�T�N;�����J$�|����W�<b�_3캍q���(�i"m�D�N'`��f��k^�˕B��c�O��]���rr���5p�z�s�^��=�{�v�:p���"%.��&���Ȋò��jE���o~�)�!F��ټ���9�0_��W(��u.!Z������ _�&���@�5�5:}1����COa���KD�5�l�����o�6�)�h�r��.g�Wǎ�B�ן����-6x�&2�(.� "N��h�^b?)Иly {�$�c�5�>$NC�����ǛC3��9g��B��zN-���2�O��s4l(g7pIV��/��E�M���-L�
�'vΚP���6�$݆�1�=Fz!|�̤��@&��AgU�	��KR�3�V���:2ǯ�=�-o���\h�C�������bR�8&L���e*'�퀼��������l,#'�[�h�R�G#U&QQ���r�F��i�|H9!�����t�������"ʭQn�uz��@��RS/#�h��Q۲����Lp{ج�,x�k4s~���a��Rr�|�
�á���` �V����Ű�%1e�aC7C�������n��(���s�68��x^�HG���8gC!h�Z�Ҁ��g�W��+���)�M����K�d��M�Z-�o�bo	���-�{*���Ȧ�#88-��2j�-;bJL|���b�e�Gc&�;=X*�G�����kd@1�}eCL��z���Oq��";�w�a�7 �Ons=�4Hzy�e_��:G������q\�ڥ�����Oۈ�>��]IKQ��t-DU�M\�p1�#���TNG�՛�)��У���
����&�b��[}���,�����y��kn���3R"�;�3�re�-�I\�����"��k��'z��=��a��΃ӄ'������=]_MC���%�'��{d85����~�0
8���`�R��'���&±��A��p�v�x�Plh��x����iL�b7���2ૹ%�\�]�5F��W8��<�x�Y�ͯ�J��������"���5�=Ɉb�aZ��h�[�q#�ߠB#7}3�1������E*��ҝdT�J-V/�,:�WeO�7��7M���r��mO8O^&J�֘�J6����I���3nܑ�*dW���� B��B�Ӕ#�T���a�4�{�(�l���̳p��o�_��m�d��,B/u��8�$�R�o�5���ľ�� A��%�^KS ���A;�^�X]���y�ޡ,�~tu,qY�5 ���Ճ�K�l�V���(����A"���)˷�F'��aoF\[��N�r��<�[{��Q\ʵOO-���FN�D_D0_a�0D\�d1��T�$ͥijR�PGr���=�A���4�3U�sҬ4C��#->��G�Bq��;9�r�f�h��L%Pj�+@NnǑDOq@ ��Q<�I6� c�Y!og�:���Щ������:�!S4�_U
!0�Z�������`Z3P~�3>���|�3A�.8��q1��-+?:��>��Rݥ٠�Z�����JC��WRj���{F��DB|�R=����q @X����E��ҷq�m3R7�Tc��4���!�[�
^�n�?3�-���wZ��i��JR���>�@h !ŴmՓ�P�O�e$�K��ԛc��<y�*���w������� �������]n��0��h~K��Q+lס���mn�W��<� ���D���Ş��2�:�9V>�/���6���P�VҐ���se�@	�ApZ�1a]lf3ɋ[0�.�����Z�,/��1V�>��c�/���H^�XD���,ȂmA�2���[+�*�ȩz�� ٷ:�o�7K���Q^ڂ��hU׾U����"�@���r$�k������@J���cG�3����آ��քd�vh�o?��&m�n�<`K/��x��$��V2+ys�_�kY饧�C�Ag�ݗ-:���䎻�/�x�op@��3U%����$s��ad������-y��Q�߁�� EƸ�t�s����$\�8���j���\�� �|~
�iRt�7T�J���卹%uO�� V]��KI%va��b੏���\�����?�SIo�LlX� W泑IC��nTB`mꞓ�S@�!�=7�`��-Y(l��uwz,c��4pv�N�W̼��a�a�Nǟ7ڥ��Y�.Hĩ<I�nt�1>�[n��2������wR;�^@��-x]"<�*~����@<��esP��S-�x�U�T�u�F]J��ɢ.b0����1drwm[\1ۙ�撖-�&_^&.��cfb�+-K��[��_虫#}����--���&q*e.볨��`�i$��ZJ��?��8�䢾�����R뾨H�LЎR�Hi��p�/��ٽʩ~W��i������i��8,v~N�rl ma�emz����� ��di8��bd�xQU �C@��x�'���q�ϯ�pUdc�CKُals&?B����~�X�P߉LG�~KoRuU
���y�j��s�oJ��=#+xy��� �b'����2�D��K9!�!�q�+���#N��1<����Z
>7��}#~�z�]�b��e;�x?����m�ſ�f�����]9��g�AF�i��ײ���ZIK�Y�C��k�^cl�E�A�<���:���wO�G)Mǆ���|�,���7�R6Żrt��T�m0ɬ>�[[��g���Y�l�k�']=W#������?�L�zk�Rƕ]P�Пz�c��֣��a�̸\h�Z̚؄+j�u��9�����}"�zR-�g�Ծ����^fG�����Q�l��b �
Y�1;�3Pk�v��l��QK�<?d��!�4FI��F�����̪]�(���kl-ۃ�P�BG����MfC���~��*�=�҆���A����u/Z�P���U��d�d$J�kp&J�:�ꆷ��� =K�������^xO}`*d�䅮��4*��E�QJ޼���c}�����r���YܘI��p��2_l"��v��!�p�J�$]�KU<�fGT
ߵe�٠���6\��w��(�$}\��ď^��:��s?�(�ܿ�&�U�ٝ�s$0�H`�h�=1�~.������%7,g�%��R�����L��O��.�"-���
^}K��Q���:z$��ofn�tw�J!����-5�b�u:sPR	F��r�esv����t��S�[�˓�=�%�1�Z����S��A ��תY�q�t��5��*����&��D�a�K�'�ټ�ؿ�y�Z�a�<|ګB�2�7��Vƌφ,�|�&hH����s�I9S̡2UǙ��7Ϧ���l݀�]%��RF�;�")D�^�h�V&�-K�
���
.d�l��1��I�N�*lr�❖@yL?Օq5,�_5�˹����O����aY`�����B�Wd<�B���,\dr������P4l�/�E��[{y����;86����,�ZbI����=��J�W�47i����<�h�ޑd9��=N��$�ך r�4�9A���V\my��?�\L$3!!vl^���~��,}����k�u)ϛ*���;�)�;d��D
������&\C�\<�W_e�e��pfTV�Wz���>���r��`Je�l��{�t�WŴ�z��"�����������Iqo߁���'C.А�h>"
i�g��I>���[:��p�=��5��/8+0F^�c�M��Nw[_�괝��Y1�݀V�t~q$XA��W�0����1�W�	.��`�����|d*�����ɷx��t���,<Ψ�S�1<��%���+₼]��|�w�Щ�������.�-ʾy���x����8>B���m��E��۹�M���y&��F@Γ�G5�'�G�b�/�!?�cT� ދ*�hfw8whm�M矽�x�i�`�Z�r(�⟶��=�78�'�;��~nW��7H,���9`ӯ�pO�0}�Si�O�O�� ���PbUpѲ뺷��DA��?9N�=�Q��ԯ GQ+��������ZjgZ�k�38g���h2�{+�4�����"}�@#œ�c�}L`����}����;�g�3V�d~b50��7���i�F-���-�8�����& tk+�A��A[�=�p��s��ƅ�ݖr[ F�K� ���kQ6��rQ�	��|�̀aw���:�'��}������J�����ǥ�-����j؞p�O0�;�ǵ�e>ƕ���ﹱ���\���qςH��Tö
i��G"/�㾭u4B�~w�6c/f&K�d�V��l#R��(WO_��oi(8׸Ⱥ�ٲ`�'������Q]�(sWu��Ń�^[�����N��U�q)��|zj �O��&�����T�)b�:���׈^q����y�(�ϡk8��Z�"�(~���׿gQba �z^֝[�b%��� /��C�oX=�0���vT�Dx9�o^�jF~ Y,�Zq @`3����Pܑ�W�v�*��nl���=��7����i�&I��ġ��r�
�x	$�+�����Μ7��� Bs�S�F�҃J*�w������r(�E��pK�K���S%�}4^2F����o���^��P�UG9q�2e%���S��Il��-�E�!�z��m���C�u�r���S���>��P*�A�;V\�Ό�II]�#Y:+ݹ��q6��� �}M���>F��4�u�'Mz���hD�������t>T�h�	O���P����_��j����Hh�~&����4�yP���7�9���$�M迬c?�VvKvK��ys�.��(=VYR�X-��Xץ�m߿g�CuB�ș�>��~a#$�Ҧ��K�U��z��P�Ô���&��{)��6d
�5�t�:�?q<�,|�'ks����ޒ7�'�(���,^���3��OƓ����r��h/��n���A]'��2�+hS��XqQ��8���t����"V��G��
�Db`��g�b���}�P�ٯ�Ybb=|̷m�WS z��a�蠂 v�����a�b�5^������^$C�����'�� �<�G�6��>���:���k^���0J-�Kě�1��#bg��K�݊��l+	���&���~^A�a����`]���يT/�6���#y-^���x"�񎷪֨g�[���̴OpdT-�1�֭#p`���Cʧ�!­��nf�(�Ʉ�>��$p4g���y'3ޒ
�d눼�����~��6GBK�d����^G/�Z�@�7��Z�8�a8ܗ����+���Ӊy$l�_�a�nu����~~ŢP.����}�P{(V���1��xR�S�ӱ�-N��6㩏Om�kP��1���W�[^�~è07��oTÓ��10y*-l|>n�S4���s���<�ppQ�3�b�m��'J��|���;p�B�z"�	�hɳ;጑IسT4&^˾�v�d+�:�:��h!!��P�s�%OǢ�Gm�����ζ��ˆ2�p�"R�4w	�t����g�Ny~X��˻1SZ�-3G=g��i?i�}}WdP��لv"�Ȅh�^)�9iB��l�R����b�X��s�G��0��`*�2~��N�(���@�B���i�*w�1ŀ�M�2���
�9@���������0�����pr���ˉ*���`����QI�?Ub��n�3����x|�)s�AK����]d�B{���Zu��|ɫV�RN�́@l�� e2D��1d][�]l�~@-m������n Jd���w}������ա���뒍�!A���.'�qN������'����#"/N���i-�� ��P��&��sw�O6_.|�&U�t�=]���A�G�8�K~)�9�4�9��D�2v�����"Zw~kn���3)���`���/���B%+4�"2������K(wT��ip�5�醩��j�_�~��|����U�lQ���?sE�r��Y�.�1/�����+�ZÅn�v0�SF�%���E��/.��!���.��.ۙǮ��5G�:��z�Q���@+9(��vk���?6u��ɼ����
�4�Siiu�U ������)0/j^y���-N2ʅ��`E����d�1Q�0_'�t�ȝ� ��O���*���z~�,�B�����ܝ�n�a�e�~��E�sa4BH���R�:	'��w �_g����CM2�s-� ƽ�E�S�C�8����}~�7{�T?	��5���az6t�"y8��ӷ=L���~hp�HB��J)��a0ɠ;�}�����mm2� FL�����+�)�5�����Çu5տoX[��sI�pR��{_�}=��iZMbI�����
��P¡��Du�Տ}������~��Ϛ��j�'��1���}��5�+U-�}bY��a9��� ʡ\)\�o�����Zw�{Fkv1%�����c�*�	w��xt��.y�A��W�vSd�������<�tG�,E�ۯ�x���wdnq��
}���J�: ]�(uTo��j$I��7 �v���k��p�x�E�B��m�+��h����!��CG�"��$�AٜM��"[�5����]D-Xaۇs���JJ3�ޥ�eH����XyJ{�"�n�����"���
0�<ɥ긵�I>��X��=��!�U��ʮ�Rcv���/�NϹ�{���+���gR2�b��4�օ�;��vӖ#z�bDE!+�����zyhQ��i]d���X���~uZ�� x�v�\��<woIL�=ozZ�K;�]yV.�)e���ݻH�3hy��D"�,�h��R�+���ǭSTis���?@��� ��ᖏϿܯV�Fm��I%#����S��ɵ�`L�`7��,������	%��]��lV�2�~�\Y�{1���z|t����L�e쨊ᒝ�WI�I_jS�;�CO0�\��m�B��/���ް�`W��.l�ĺķX�])�\�|�gԙ�I��C<�0�!v�����K��?���V%�%�TZ 9���h�j��b�yy�����VF��쎵{�5��c���d�?���ඇ�;.�ϻ+�HI�������xeFr��Gd�p��^E�
No�h�ޯ�d_�	�ەP2ƫ5�[�v��ZL����wb�`/����rw��:	+<�/zz�����)��P���5�_�K��3�q*<ᴊ]�U�i��_��5	���y�]z�?�1�a�~4d��p�0�2�g��Sⱁ����-w�{d��GꙊ"�i�<���šI����ҋ?~#�>W\�g�M�˺&��M9�,��_O%)�p���H�X�8й���zp@�L��|<�������\�'ug��x��^zz�h��X���Ƴt�viE��^r7�$Y���8���+���(�������� $����+R�V���_ѻ��q�W��<tbO��~'�/ ����T�`��X�����#]ٴAC���q#(A�̺^��HGǱ6׭ފ�ˉ7l�#ZJ��DWE�k�3���
�x�q�T�px ������O��d�j�럹�� �,��'���/��ʁX�c����΍�@���h���=Z�ܽv�>j�w�p蟟��h�=;���2�ؖ���Σ�\�4�_�~��MS��D35�өi��3�%+��/J�.�U�Y#/�gO|O�P=cbK"1u�s�������(�
(�6�}���ɡ?�£'��j�x�sV~�%��a)�u��h���f�	FQ1Mc��P�y�U6�#�7���jud�~�$;9boI1�f���{I7�X��-!�3�3�I7L+�q�U$���#�ǔ�9H��Y�g?(^9o>b�{`�8��'P$�^�~�^^&���vD��� �	i�)����C98鐢��ټ���{��d)������~Q����p�퉰����*�3�>�q��8 �%��@��}Q��|�97d(lr�ۣ��V�#*]��ǪObV��HP�%>f��6��g���lW�K��C�E����6�@����t }�5H	d�����>R3"��Hm��Z%�;t���=�S��%$Bӑ�����u_*ݦ���]�dL'w��mP�,�m^�uu��bS;�-z��.���Z�S�%d�h%":�m���&�6!�W�k�r�7�߬]� Ci+u�ݸ��-UGQ��i̿���V��)�ˣ�9H�t�����i	..�����$� ���<�����h��ΰ0bH����.���.�5F�qG�s���CG_��YTh�4<CEm�G�q%4�wX-D�'SN-j�\l��@�'J������]sv,�l� Y���괛��_��G�yȴ�B��LIp�\k-H�'[�BOM��_i��Zg��6ߔzm�RK�q��bn�KD��.E�����+����
��\|>q7s������+���2Z�s!�l�2,1>� \6&�}�G�;�����=�{�;�NQ�]s{�~O�#�q�ʁ=��rH���g�v�[�1����9�]
���	�5O���zF����N�C)~��f�Tq��Q��I-}u��R�Jǲ����aN�D*؃mBh~tFZτ�'����������˿�TܼLq�>;�dl
����jO_��75���^�?@؜�E*jYJ�)���DA�Km����E&�!�
���I�h6g��cwr�{0�E�<�S�Kn��=��v�ʴ��7����-�@����߆W�X���ِ�F�0� rd9�6�,��/�'��K��h��X
-,��ҭ�!��Ք�tA_��=0l��kL�b�/(���	��[�_�f���+yZ��Q�'����)i���}�y8��zQk����/����"��݈©��AK_�*+��/����U��W�A�D/ѵ����aGu����0��O��Y���2h{��#aMW	_�P޾ ��&�i9M؞�����+�b�=E��qc���ګqp��`�ܿ@UW��`���&[g�J?liS:��/�47x�m^؂�	��!+�:��*<��;�;�jJV���|�: �۷T��/�^�R�5�5�s��m���]���BrqG��O<��'��!��/ϲa3��Q��g�I���A���Wv"L�
4��Ccό��(zFם��/��;���L��q�(��Lb���+^�w�aP]S���ɂ/��׉�`�1s��Zw��4+�!�]�&��<����x+W�5����>�[۹pL2R��O�llA�X�Q�3k�k 9�l�#�K�S�e`���`)必�]� Y�}?���Q��a��1a��,�T����z6l���+�PGt9�,�P��%����+Xɳ��s���Y�1�2��酤%�r�������5��������Z̈́�׀��sv-&�T�nԭ��\^CaZ���	�狣BoR^���r[��*�`Wq�.�9���g�~���X$?#���3ю ��Çd��9`\ B�ҼqI���L�I��Քj����@�o�&�_��u���ְ�ݭD�j�����d��+�G�Z�9;�㰾�d���J 6Z��upXƂ?�#��1�4+��fun�\W����vh0��x��}P�{�O�>���V��J8)t��?�KFj�����+��]�׌�Н�o��͏CeӡM������jS�Kc���^�{�'��兡�˸&Z=�yL��^)����gQ��o^�����4�N^mS��x�<Q<?�*�b��]�6�5�.�$����5�1�����:�Ԁ��6�#���Z��i��!�*tߌ0 RGM���/����w���vtd�-W��>�[�YQ�m��t����3,z�FB�Z���Ǆ��0B�!{Kl;	ﻦ�q٤��u,.&.k-�'�x���e[�\�s�zm�H+���I��ݙm��[T�1d���ֶD�w�z��(��:i�a���0�@`�(խ����������aTv�l5\�m ׏o)�ǯQ�����,�[tJp���
s!��&�f�WX�]#�,/�D#<!¬�����Y�%���f�Z	�H5� -�ߔ��G�B�X�$+��u1�O��� �E$=�������Z�67��[�����B����0�=,����{[���J���w�3�=D��
/�:�(�)�Q�5<}A�I�D�"y}�M꒭�'�g�w�t��̮ǐtQ/�+j,|�=o��#k����ù
wB��]�G�]�͛�% j�	zA�� |;�*�0��k�&�Z.�z9dm'���ҋ�m!k'��e��� ���a�����M�w��Ș!���A�$�m�5�agQ�rP��_�zgo4!�Q	�  ���>=���#H�����&���b�;w��.�e��<��
�ե�~NY^�&�O��-�bx�W�������2 ������y(�y��&��b�����t
���z��i�j ۭ5�֌@!�M==it�Ǫ#����8�o����)����u��>Pέ�p�Ho��:��9�+�9�L����&�fX�.�����YgI��!��<^�&UG6mw����*p�v����U���@��o�lh�y�z�G���ߣ�-=��S��rfq��}L|�e�v�3S��.^����"��5���ZN�K`��Tw�9�A>A��m�h�"չtaOx-1��Х/fB^�eY�����4:�����$�-������#h�)G�g:rlH+�m�w&G?�XWi&�c���x����*�x�/��K�$x\K{�4��F�`R�s��0���������N�?їԂת�{}��9t�����H��Bo�U�wy\��~qs�Dqٷ�������U1i�7��l'�c$����n�#0�YvE���>�����������^(z-�~�έ�"���s�ZeL��"ƺ��;���m�Z�Z�9�a��� Y�x)���c�:4��	����l^�n�"���:U��v�|�XX�&��E�m���C̽R��V�jv3��փ��] �_'���I��T���l����z9M ŵ��T�)z���9d\9�g��v+��I����#W�K��i��wv@�b�I g��P���P`TA ���Yc6��N/[�D��_�Hlw9�y��]��Jj�G������ȓ���
�n���5��_]����z����_������ 8�� �,�sտ�	��X����ʗ�'��C�ք�qMjKɕ�VuBQ;�W2]�����!-8��#>������<�'�q��g�T*7P�����Ŋ��3�����FʜƌX��{��y4��ǊH�Ғr��| q�8ǩ���r���sݡ?�_���ۑt���-�����m�e
ŗUQBE�Gw�P"�����s��:NW�0���F��9���T)�a���2{� R����/k�T��Lz"I\i&*7�(9".6@�Ǉ�Kg���XW�1I�:�l�K��{X��'A��o8w@4՜�e�y��XR�`m.�frJ3X���A�O��%
P��"��?w)A}j�y>��l=�R��l��s�G�4��;T�zCT@��	�̄��s�MF���EM�o1\�7J>�d���n (G�����+��+��7u?��C�ʀ}��N���Q��H�_vvD4�C��֌{�hS~���F��w��c1]��E�H87��R�o��K5Km�l��CK�9	�w`��_�����,�4z�o4)��Z��'�χ�@n��פL�z-B��)B����KP�8I-��"ϱ�5�nXާ
��ͼ�X���y	������>�>2l����#�U+$϶����B��Y�F��-�kY��A�w��0"���ď�9��6+cu���k{C�j�R�Ox��/�
���.le��C\=(�����V��� 0��}�|qb�͕����޻�$ؼS��$��	n+m;��e^>E��+��q][Ϣ�eH����c-|�%6�TN��-i����3����9�S�s��]s�Xr�p�9��c�5�P��z����?�AZ�o~������nSƅ�J�:n�K!��E�p�g��z{�D�e{�gJ�y*ۋ�{�2�_ŉ_b����@u��g����8�c����H/�g�<�uǧ�ª��H��{9����V��z[s�P r7��d�D����ݬ!�`�ܒ�s��Y�2�M�������e���Rd-%`xV��3�qH�4�r���TҠ.bq��ΗK9�*��v��&Y �Q,j��=0�=J�"HI�������V�:�d}���㓤A��W�K� ���Z��>�'i�+�e���A9�Q,Z�a��-1�ڨ���A�M�؏����N?^qW5Y**�4��B�}|rW�BqAfvA�����^u��6�'O$7���o��X�V�%�~;2����Pd�� ��.�j,h!�.l����	���'�ت��j�Uca��bN �2;�hȧ��QZ� ��p'l	=}�6qD��p�Y�~��o &�O;���tuZT�=ZE#-!))��!V ���3��Y��"�&��z�nGy�28�1�uT�~k��;��j�����+����T�����Kx�]7����#Ivp�5Ǘ�CX��S`�d���x�t�ݜ����߾��a8C��fh6�Ȼs����f�R��J���(�T3wW@�� d�W�wGŧ)1[`�|�Z�g�� ���2��}1Ճ�����ٵ����eW{ k3=�^(�W����wtBę)c��A:�'-v��W����1ĕ��ȳkɯ��ӫu���̰���Nr�x�F���}��,��B��$�=#�zq��I�b`�YM�AL�����{���6�`wv��B�!�rI3l�n�#�$�k�^
������H����:��vĘ�����QZ3Du�@���Ei:����#_U�� T̅���[�n�	�&б���žT���~2==)G!fq��g�E9KL�;b+q)�Ц�y��^��}q�ų˖�(���ҽ�(�6����B�,'�H��)
b^�T޺8X3����ܦ�_���
�N" -�QtEd�5�z�P=4f��V4ǈߍ�s� (|i�>?�[�y����b��d���ZE�"�<������ŷ���j����m�+-�7e2I\wd{��!}Xo$��l����_�_��8���hxݺ�2����^F΁�CXF�5/�f���xA�eL��,�u��rF��n�id�c#��xY�KTdQo_v���������f䌩0�&pg~&F<l9�Uz� y���nI�jA\��Pћ)	m�6�ڣ[�ֵ	���q>�'�b
B��X@�v��Ej� \���>������V|�P���b�<*�(60C�n����]�㜭�;�o�_�v��
�ԡ��u!I��ę��c,GJ� {����}W�jN��{�XO��j���� _���ِr�
"ÖUD;�}��*��=%�A箽�au�<Fu�D�dƱ���8���%^%~4�n���-�Ѹ�坩��x���hԐ���}�����l*W�?��5�M�ʙ���O0�Q�������z���IZU5̞9;��g�[�L�n�J�1��7j6�%]ek�ydD�"�)_R�j��SH���L���+m�J��=J)V�n�V���y���La;��tQP6Vv2���'�����Y�B(� Pz���w��[���2��&i%�dY2�)A��Q�2o,�*�t�\�M�2U.�-b5u� D�^d卫�`A��*co|���R��w�J} �RЁ�Z��B�I8m_�Dm\���ZyS�|Ml+e�������ط��,������|8�32���m��߬>�y�i~q���8�=Z��x���:�<}�t"��Q�h���}��;~�8�S��0c���c�v��������6L��{�əb�cݬa�%c���/���fё	���:�˳ٚվ%-&�:��U5g2�e�d����DR�c,��ڞĔ
I!3ͱUL/�*�M+j�� D����Gt�?��v��::��G���	|&(t� �w�J ĕk��>4	2+�^�U���W���4Tj�L$<^�#����o	&`X��y���?�7�{^u��	OY\��ԧ���L������^�d�z<v�G%�
�T��2�N�&�Z49��Pڧ	��7!�F@����\z+��+00��@�o�_;̗����[H����5�#rx��V�QŜ'��'_�#,���$���� �^�Mo�m?�',��u�+�-�Ε�G�~O�3�cߝ�H��s�&�r%.�<�л�&�X�6�Hք<��.<�D�n�3�]��B�)�rF�lpȡ�+��l��v,�g�)�o)5��-��
�V�	沣���u�c�$ZɈ�_s&���{!�̀��o�1��	�^�6K�Y
<mC�v��6����7y��Tlտ�Һ�(���uw���#	s:"�:t���Ƭ9h�����x�>�� 4!]��o�V���iIL���P'Ȍ3�3P�%�~8H�˘���q��kI<�n�2�Bk�\�%���tCR��a{}bS��3&���&���s��
vU��>�w�{�p�:ص�L$i��Uu�j*/��.������O\��r2q�Xp%ͪ82���h=!��c
6t|_y���?��	D��yDB�Ĥ����������1�j>l�t3�c��^҈��$��\8���mHy���{/�׽������]#3(jt���,�DqN�L��Ň=^��@��쬁��h|	����42^u�g�TL~�z1WF"L�^<�dA��9�
��Y�#&���Ie���s��y%�E�
�*�e�<�ż��5�s9��!봛Hwt�^�l,?T��p�>��PG���u�x����:��g���@I�&4ϙe���������
���v�r�g�����U�?�n���H7jH2�4%���ϲߴ��[ QuU5L��:w1�����D�3�Ge.�i�-N��&X,�M\s?R�\/�p�o1�א`���#@7]�3ؖ�?JB�ℕ��[�Ǣ��E%��M`��|�)'>_�b"���m��zC��ƗqiS���U���s�k���w B����l�+�y<>�+;��5�tI�� �J�0ږ�f������7�c�O)��Ǔ�lb��0���"]�sV�Vٓ�Ɵ���ـ�Q�~�:I�PWWy��v�q�����n���9��o'����\���-Z���t����+�?��V�>%�$��Jy��E�ĩ*9�k��~�`Y�Ku,0lT��X}�v��2`m���<%$ee���ٰ|��5��B�/��~�IgP�2ţn��K����_��eJr}��2��'���b�&v]��M� @�����C��n����ֳ>Y8�6b��z[�Q�y",`�_T�W<��I����t|څri�l��ΰ�ھH5�K4�"7@�/ĿvC�ti�Y��{\~��4�Fx��8*qG��hi1S��%Rv!|��/��t0׫_�.Vb+�$[z�)=�@m���~��)����c�#o�%�lc���na����]^���k,b��(�E%}��,h廹���W�V�K���p0�\
��=����qu�\�_��%�|�#��L:^�;-6�o��8��+�1��U����牸�9��^����5�0�"����� ��-�^{2�<���5�
��z���ξ�u���vl��,n!G	�ӈ�<��!��n�,���[�g��8�f_����TUWO׎`9��o,|;U�!��\c{C��W����4&����n ���Ĭ��L��.��7Dw4gm�J��HH�V��geշғ�} bۗ��`��ZsqD+��B��'�vh��'��56��e=s�cb�L����xP��k@h6�<[L�E�C?��T��Eh��I�?�o���gY�0�(�%X�a�=]\F�]j�F55�v�c{�*�7�+�v��'���l]q4k����� |������R[�,�D_��&���%-���C�� sT�h3n��)�����}y�nIK���mw���U�|��^��1�A���z^4��e��C��nRN��K�w���Y^�.�tؘ8KJ�?#�0���~C����> �3$=���DM��PG��n��!x���WFfɏ*gm�o���ГK��h�vؾ	E��%��ŁE?���P�Wu�ЋPw���E��G�F�G�cD)n������������=�?Q7�_#��n"��a�m�eNɱ+L�Ԩ�	[+M���|�߈�1�Y��>�!�4��vxԤGP��>�y�.�����.�:[�r4+�6n����$���X���A�.G��i�kiǶ9")���\(	?� s��)(�$4*X�C�uN��=�I�ݜ+�S*�O�y6�"�J�%�ฃ�D��pR�m�#�l~A!]��R�4�6ڴI��f�Z:��x'b[���Oϛ$ ��T�ș�k�&"`�&��gޏ��=�F��92�*��Mx!Jr�&Y��ԜN�3��j}�@�	��Q���6��+�� ᧍�d���!�[jO1ΰKV(5"�X�A�D��ň{Vx�j./�kf��3
�uM�����j���B3��e��[N�B/�S��b_9�A��q�1_m;[�Ӎ��ۣiJ�&]�DH���y��qR?���7�,��*���$h��9�	R�#��_�0f���j��D7��I�-�l�e�n��}��0�T'�%�Sֽ1��4�-�?ev���Ae��u�x�!��[�zs�+>
�h�՝��#�"��8���U'�B�/<�\;=�(��R�@��M�PXcv��'�q�<鯂p­E�������kq%Ɠ�ye����,���T/5�j ��<)i�f�Yi%/2�I�<�k�[�]C<^7�P
�Q,����	 �f�����q�{�;�`��7z�0z�[ֆZ�s�rj2S/��f�P`r� T�h���P�^k��J�P�SD&=��V�	ȫ���{",Ii�i8'��R�}���f6��ty�8�
��Ա�e���t�pg�8� ���bҏ�!iw+����k�����y�z�1�v�F,��̈0J�h�)�[��(�C�w�<�� "H՜4��E������M��y�=�*�ۙG�ғ�Q�5�W��A������r��	�����~���8�3�VΗ�%9�D�= �Z�{�p�$MɂdOV��s�̸����\-���Wĳ�,l=x����H�v�$q=d� W�CDѭs�Fi�VO��4_L�<1V�D:E��U���.�(2�,����3�t�V&����w$�W�7L�N�|����m�0}����q&x[�i��F���B���N�2iK)�u�@L��9��;D4�-~����~��s!���`&�f,w����%�JI�[�M�%^G�Jq�?�_��&fI�����G�G~8�ی����K���� ,�ĝ�R�B7���������Zְ�³�����+"Pw (W�&�$��Y*��e4|��f���V�j�4�!&R� S�Ҽ�EFQ�݋�b��j5�y���C�7�s�'48��< ��w�E]("'_�]"�qa��͡�H�;�;��m��!��ڥEʅ���#��ǝ�x�~�
�W��	u����?%���R5D��
���ˀ�@(�78��������m��L��w��
���.����C��6<�Nī�z������J�7m/��p��E��LO���8Ռ#T�R��~���E���q�{f
��ki���&��j�B�_��Rב�5)x�ܣ�0`�ƾ�V�X�������~���[0�����������x��!U��c�4�l�Z�KD'	��|1�����1oTE��W�������Fb�Ci���<�@Z6
� �/��QX�-Ċ#|G�ۄ��S�jqxj�5E��wn�%ˡC7�n�P�&~�*�,����ni��}r�3/ �~��m�/W��Um�2�]�Q�8!�(8�Y6"�Q3�u�`�#;kϖ����<�6�d�l�����6��:k�U���Q���GT�jd���d���"1�DY���74������7/���RBx� D�#�Z�XX�#�����NA�0�w8���z;Z���-��k!n�}rMl�m�|`7Pu*�8�/����qL���M�]�p	�_|w�
�0zy����I��������kк�ES�ߚS�����Z���R�O䬺�Y�E%�3�PI����z�"�7!�<Bkt`��5O�%v�%��I�x=�r�8���NX!����p=KV�I�`�*Tܐ�����Qb!޾�[t�5y�jG�c�Uxe������e��ô�͂��/8�	�.��d��#��$������!��	��9'&�ƀ���iɡ�T\U%ès�Oi�f��>�eS ����3ȩ�S�<���V�e��:fu� ��������$kӎ3�~!�6�,��vq{�~���͞q�1�F�����H9xQM���0�~9��}��|/c����&Ul;��Zu��x�]J��l2ۄ2f�SE\}\���.��z�R���m�]�sAh��F��{�H"A���Y赒X���|΀8�D�$��uG��,���UW�Sک����-�,��kw��#Ѕ��Ԣ�&��p����@V��
3Rg���E��������WgР�G�U���Mx��C�$1�*�Rb�� �=�C�a�4�R���j�їN6b2�͞��v��@��f���l(c���d�jPBȘ�gĚo�s�n	�NS�ǩ�|ն�ּ���ɛ=�8b(whM�&Wo�b���xJ��b��=T; bq��Qc�.oe�`���Y����}������{�]����坻	&[�,P� /Y�D�N(eu���*���4�ފ/��Vs	��\p�*  �g �q��9�\X,�*��D� z^P5���^=a�S���������@ڗ���I��uɥ��ϗ�`�S�0	�uR_[7����l����3ڞ8p�O�(N"*�1˷�5�����1�r��� $��d�	���w�]w�D~������֭���#�(�]{f�!���br��K�E�T����=�l�7�AĀG�����gds���y]1m��@KQ�>�(���ɟ�a�l�l��cX�C��ؠ��Ʈ�t�#p�A���3Ֆ	�C�v���b^lD��!;�Ţ`YK~�z�$-���q
�����E|ot��Ȣ�����=g��o��Y{6��\��|��'XzZ?���u�cYX8O>���%+I�`��ئ�ۓل�ܰҰf�0
�B:�
�6Y��@��Y��P`c�u��ܮ�0ww�w��:�f��^�C*�\?���p�K����kt���SHB",F?�u�J*1�����������HON�=?Eĥ���C��%���� ,��:�} ��͵=�T�[���� 4bL�ju;��v}04]Y��T(�BHsi�S9���&�m�$ӈCΦk��k����1��U�[��'J�F;"��;��ݐY�كj�W�����P�Φ3���Z0�(��l{ŋ���5�ˠ�)(�~K�M��T�q�@L;G宲�����r`�b�ݨ�{f�� ��dՉG�*�s��Aq�e��T{��i��]B�����56��o�b"�z)!;�7\Fp:-tn|����ݫ'�{oq����x�b��*���∢|]��+�m���#�ɨ�q�����2�1�3c���½�n�±�](���Ǜs�]ȝ��/z{n	�tMA��?t���ܒ &ιY�d�pXԂ/�]n��av4�I0�n���GPqNf�略#bO��f��LR/����T`5!��0�I�W,|<
�+t>I��R��-�Le)�:�!!�y����f��y���b�ɧǫ�s�sT���_��/������$����RO�kkj�F�'��:Ȁy�5��X�(�i6��ӹYG�#dk�yŝ�s�w0ef��� �1F������I�L�u+��_�l�^�/�7�\�����"D����As˺{��|�Xi+��3��a����WY��h�}$��7�F(2Y!�>���wx��Z`�߫�Ut7��w�dغ&��#4Uwp��IAe��� 1�X��'z�b)5|��;�I���q��d��}\���������1�<f��=��irn���mς���t�����;�1u-��Za.#��Q(]p@f��I��2�e��2�k�@Q�'j&+�2������O4��[�sel�0p[�L���8w"*P�%��,�d��m�)���3f�췡ơ|�w���?�S`�}ݳg[L�:��i��|� e-I�e��+�����9�W�=�2 rf,ӿ� 
y��-0R�{���1x)ǅ6|��0p�,�I��fh� f� ���t{y��^1�3�G��0��#�k���:g�=����\<���wё�B���f�~��Kk���+�ЀW��i���FI�]� ��6A㈾�/��?$6QtL��f0�L��i$�Aִ�D L�xa�7��'��y>߭������Bp�{Բ�G��_Z�����D����Z���S{�B���!���P� 5��yNK8�I�3lٚ���Cgٽ� �	VJ4#��~���8|q�ߟpD�
�qqђ���2ܦ�̉�\ZBhR�e���L���\����0�� 夜� ���u�q9�����7'���R#{�ܷ�'J�_y>ج��W0.�נ o��->�9����Ra�`4ۡ���IZ,*O�"��ꫥ��4��i7����@K���5璴X-yW��@ry��ᏺB�wv�w�f[�(�8G��Mm����8�e��/K_�&��.�őAG�X����Tx���r�NV۩�����u>�y��̼��#�SZ�
*"����$m\���y:�v�͞����t����z����qQf)d^R{�>��x�{���/��)��o;(��>��[�jق�tQ��	o�;�w��;-��N}��(�r��d���+��EJqfLM�8��y$g�.��¾%˟�&�S(��n���+��"<IdpCZ�Z���|�k�߲��X"˰�3Xa�e4�7��B�莈o�(��qץ������p�@���D3�f:����d��ؑ�G�@����h�-��:��$���V@_}a����ƚm�����-Ŏ��H̃'��٥��L�l5rmD���v�j�X���!�6Z�*4�Q��������T,�
k3������2��9�o}3g/!2y���h�pm�����I٥T���L��ƺjDZX��z&TQ[�.��cB�+
�$�6�'�!��%=Ŗ'���.��UH�4��Z�;�$5*��`��d��(rԥ�Y�j���6�M�.��p�h�ޏǬ�b@��x}��Ht�d�Ee�@�����m�����p6�ґv2:D���G�yԜ�M;Ŀ>�Q{W�U�l�z�V�_��7il#�K�:�!��)��%%���3�e�]:"b�b'�z`4�~OU��5��-I��M���؍U�T|�w�X&���.�����<,��D��^q׎'̌�l޴0rQ�=<䦘9���m��b�}�j���Ӝ�z�A�a?\��M�.�׽��xx䰹#�ǒ�9"�!��a��֑61z�
T�JR[�)U��>�T�^�N8c�C~/R��y)�k�B�p�@���-�@by��4�͘�na�v��V�z�2��?!���"�1a9��)ba[�r5B �����x�ȴ6��S�;]1*���	����wB'���G��Bg{�Vi&�?�j����w���2�S��DS�pa;_��\NH~��_�T.	{�k!J}�M�����!}�+��bv).��RP��x���p��O%핢o+w�-Jo�y]�E��'�����{�i����)��Dx-lV�i���I����������� ��Cf�s�Tg+����7�k�,��4W��,}����FNq�y�[���S�xv|�o-Aau��e%3�C����/GZ��ЮQ��%[��������)F���:�g6ڍ�؃=�w6T�9:b����b���I�HI�y �V�y�׉���L�N�0�r����iv�o�0�H MDT����~G8��Sse�5�Y�$3�;��"}���9�E��p��Q��)��i���AUF���5��r��LM
	G^��LB"|��Rزt��K0�/	U~�H��0��q��u�M����%÷�іS;���Ns=z���������r�tP��t|��OVU���7�H�4��)���Z��1�����%]<j����l6:N3�AG2�!��?��J\P�12y��t��Bұ{@�'�a�����_8L��,�'��xoR�;�\�>�n�qru�U����g�8�KrI�о��<3���4�oS�4�y]��˄?�ղD��d��ź�,�|o��)�Bz�m��u�"f��~���i�^��>��7ʆk���T����kD��֙l ��q>k^�k\x�6��N�l��|�O?4�0�9�M�C�Lي��b�w�7L�ax\�\;��M�."��׎t�j��x	���m��2����̢oA`NZ�� ��_�P_�7�_�] �ĮCy���6F�#�z�3��{j���cM�26��7��W�4��-�z�G�`#�1�X�Yt~�D��{��%�do���kWw=�O�Ѹ�k <o�$˷1A�&p8�z�n��I@��{@���(��x��.?K�R�c3�G1~Y�̯�3PG��N����gn. 96
}�zI-p_��WP���|�Z����y�#W���#�1="�~�<?�/pL�K�\��O�P��>��/�[�}Y��Y����R��LI�������ߓ7c
��U��ѯ(���E3%�t����{k;U��gw�K�_Lp���X�~�j�K���>��Q'	\�܈x�J\��S�g(��E�������q��q��0�����;wf��u��7
�ۊ�$���'��w���	}	��+��>��6K�!�8Z"f�QQ
&�Ⱦ+��=�0*UTY{��TW#����c�_s�|>��5l�HѰ"y�Q��[u�G�j�M��p��m�h��$�L
G��ݹ.��f_�3H�e��AX�h{��t	��\ Pg
�L��n�Ŭ����
���g��u5���Y%CI:�9/�*�~�e�O0($0B�dՂN��Igq�ܱ�m���R�C��6�_�s�o�p4�p�"Qf��T�/���~�	dĂ"�}E{I�Tc#=��eǓ�������Ǥ>H�7��OC��VX�m� M>k$������~>�Jj{�m�ǯ"+;P�]��9t��=�����9i�o�8��7Rf� ��/��H�2���.�pY4���an�z��u�"�bKT�k�o�_���#M
bp�h��1�>���{�?��A>�m[� ��@ ��_z��-C�-��/}��[4D8����=�'�7^������]�3�j���ޜ`�Ȕo���hUpշ��� �Y^����g��"�nZȪ>��c���(�+��°��V���o7�W��xl�b��������;1�o��gV4�%݈�1���K��R�Ϗ/a1}�Eܣ��'�aAۮ�w��VQ�w��n��'�1��Q5���S��^��ذ}_/������R�>��k���Cv�H7�O6��%����*^.~3�D���P"�H���E;�|l���$q��z���˘X�\!H����$}���}��T���NL�����h~�c��Sʏ���s�?��3pH�L-��8Za�G��᜶��0��${	���:!B}|Lo<[�;�O�&�	Ҳ�k�)Tb4�$6�:��Pk��}î��>D�k�ֻ��i����<������f���I0)���)qV�sw�� q��RP�vB|Y�36M�%Ũ�� ���)=7�:K��FX�|5?�&��%�pC񇗭��t����({�mո(���>�@�����\�э�9�}�W6N9��):ΐ<?a(�uB��OJw�f�g�$[I#�(�VG�靨n7���r���*��6�'&�EY���7��E~m�:ؾ�)��G`&� �� �"{-/)��@�f]>E��Gv>��U��c4}3a��eb��ȡ2Q�oo�`RDMd'y;��5��� �|D�/=H�e����5JW���5����n&9��X�YQ7G땧�cYAATL8�>Q
��ѓ���y-��c������;j�Z�"�a�&##��I�i�u�;����}t<�TЭ{��t�Ո�-�-��aK&L��Z׈�_�����>a�l�@��!_A���Wy����(ݪ�t@n�2y �b����
��mn�(���x�ht��ƚ/���C���P!�NU��w�8:���BO�	e����p{�`ݩF�����\�fg�����T.k_�]I�Z$K��ڴ�ݘ�����>1�|��A+o�U~˧�����E�Cc�(WU��]�&����U�_�ܢg��?j�D�z��w�3A^9q�.��B�r�p7*8��k�<�%�	"��t�D���5"�s�w ��%5�4i����� ��MG�����1�8)Q^�S��.,kՅӪ�76�A?��V[�`zo�9����D��8�_�L�-�F8�W�*k�%� �I��0!չCr��mx=����맙�vu�*J��iO��  <�v_����6"Ӑ�I*1�c�ne� `�?^P+�W
��,fԙ̢	���66�Z��2���i���:E����o\��MgE�I�N`62�Q�o[��#�����3ay����CA;��N�@2`��G&��1��Wh��ZRAG�B�,�]�ۇx���g�:�H�M	�0��&�S�ֲ�s0,���"3Z��_�"�@؉9��?xh�;�Ʊ��P)������7Y�ռ��z`���
ED��U���H���Խz��|5���Α��3Wx����U�jG%T��3��;�����ȽZ�a���>�a/t�@�i��(��C�G�]1
��ơ!���H܇��fM�@�B��X�d��<����_y䒇'>;����p�|l^����|�;E+&�a�VN�#Z�O�ۋ�3An�M[�W_W��{N��/ј���v���!��<ԡ+�]�=�g!`�tv�A�V��1$��"�S��vW;�W�T�C��Q

E��|���Zض�qm��-k_��L8yǅ��va�xg���n��3ƶ��?�
��ߺ\�l�>�h�JZ��Y��),U_��s0������FK��Ǭғ}M���-���?�0+�.���ȧI��&Tp���]�ä���p^@�p(|����YK��I�p��8b%���K܏q�S�`D/ռI�l���`���uqET"�Ȋ_R�Z�UK�~?XݗE\���s�P� ��d�{� =J���[EH�&~m,w�4�T��n6O����K�M�/���� ����	�!)��/�7�Gg��H �Lă���N�Mm38�<`�?����d��n�i��(9���˻�m�ѝ4����65Ư^{�D��I�|�K?өY咔�A��X;Q�G�ʃ��Ț��=�8.��Yvx`'���`L�� 8Cש[<��܉�&|և"�0[F��d�����h�C��
�i�D��ɟ����+
�M"j�P�,���t+��r�>���qn����0f�/O*U=R|��E�>��)��S���ګn��3��>h�o��揚������-�����`��l���\^&k�+u"!R����]���=ji��2x��-ꠕ�� �
��|]櫜�B�+8������@=�8]�OY��sr6�N�\�ߴ ���Jշ��r�u��9��@h��YF8{x렄�p>��~`= )>#&��߽��{:�6��#���4�߇�Y㗆��I�Y�*�����ȗ%�U���^7��/$����߻��J%8����T%�<��۸qދ1���x�!��h�hKC��c�s�ƚ�AC�t��$a�� �}��k	����2c<
]�6 �:�'���K��Nq}8� K��ݧ>+��7��]�>�A��,�}�t���3}yG�(���6���7N�/� W���������T|�<�"�gي�U{��9�Z	�֞��IX;7J��&P�����AUV�} �'ר�3�>��r1�_<]B�T�>y�ǀ����=�:U�:7ӎ3�m�����.�P�Ǡ9K�=i>��m�ab=����|���W��$��aqm�(�m:8��f�������~;ߩ�nTD��EI.+e�k79~M���)�(k�I�Ǝ�=�jQF����O�uU5ش����*˻(m*�:�yH�
Y	yoټ�\�	�t��E�{��)�`e�w>!l���k��0��ʲc� X.�i�K����M�\d�`�|��#o�A%O��y]73��s�td"�HHKa�|��A���1vԭ�x����rX��kPXK�	��k>�༖ᚷ�p�{�C�J��q�K��c�.ë��T�|��&Ъ��nc0�a.,w#����(J8q��v�Y(�X�4���~{/�E�r��sQ��ϢH#��ZWL�aP��'l��|ԥnh�Xr��( X1=�b6��ɩM��u�4�����%L�{x��b:w�E��25��v�{(�Tm�c`A�6�]����W8W�o�'�WG_A-�J-h��1䎸�p����*��;!����i��7UZ�`ϡ��R'Yd��Ǚ�tY�?f�������׼Q��ߙLI!���[e����d~N/;t����痗�G�SG���*��ٔ�]24o�v�Ptre����������b52���g� �}��V>[�q���:@Y�hY�/i�T	/ 55��^�ђ����*����k����1�5���Tz*Ľ�ﶥ̖qH�n�MϾ����Q�|'Y�Gm��j���u9���\��*��b��ZvAeD�P�^E�=ez�Ĕ�Z6U��C2j�O� (V]:K�����6��5})�VB7(��CS�O�Q�Y�-����/�ҍ��#�f�:��㒂�c����>�t9��r��	�xyL|�9G���V�>�!t6�P�p����\%1���L,W�&���؋v�v�%��G�nY��I�v$(��;r�t���G�[�&��a��.R��z�z6|�ESRg�~>'#�V�r�<�UkK�*�8�'��Y�r��w�4��h�w�	���o#b�}��U6�ǳ[�ݖ}�R���cʜD'��'�ʹ+�{�?���^l�h:`d��&P]Y�i���Y�Ye�L~���s���%�>L�8xm^q��L��?:bR���OԿ��ZD��k�<}
����7���pg�MRAvz����S�p�k�����r:Q�_��H�x�Q�.k�`�m�V���v(�>��I��/�<����ԍ�������2+��~��Dw9���}A34�%��W�4�v�If^J�m(�W^&؏8�#H
��K����*Q��MGr�[n;!X'��YV�M��Bw1O�Z_��ǃ[��QO�?Q�?�k>\��t��p�D/������>�b�]�?C`��0��K�.o�2��?
�][(?ݲ�}/�6��u��݄JJ�:պє}���{���+
P