��/  �&!�q]���7�.�[=Q��b
K���t�b����~��LR��j=J|��o�F\��td�c���Io�͠Ͻ��[1ܰ��[#߃F�?	���v`3ؚ�/��j��:mZ`LMUX�X�� 3,��G=������ ������6��i^�c�%�Am��^��<�J���6�����֕��**�4�`74$�xe�#]4��2��~�yZĊdha�/j���}c�O<��Ц���]�4ݷ���ۯ���+��
�G�Onx��S �����n��]����)u8���D��)X�%$�)�Z�	��/k� 7�m.��@l�9���݂�+�O�8��e��H�X��<(ᓪ������WSjl�?�(q����?�R�qiк菟�@ҵs���$(�j����n�хLB�f�Y|2�+��5L�S��Z��a�~�I�)�8��I9���%�^����]ک����v��ש�b%�����!��fs'C�ό�L{+��f��_i\��΍FC'���W{)�5S�s�_Ex�K�N��g��LU��"�H˳R
������d'!�_}Fz`\)l�6�-���h��{�yH,������:�>K2�sFV+�|�Q-��f�)��[��6sO�(�!���B�,�#���V�%foK���-���<]o�v{Yi�ͽު�cp���S!���p�f�݉��w�@��J�.+a��pK���'���Q���<XV�������w���Z�w�"�O�| �*P.^o�=z��ڧb��i�;��f�k� ���@��"z��℞�c�W<�li����`��r���Ť��y$�h�z�KD3�)4kn�L4�[�TF�����vt��І㮨YH�(6�D��_	��*I������J<E��4��"G{ڝZ��[*8�k])Tvz��X�m�j�WSP��D��� K_�n�o�Pi=����|[�6�y����[
�-L~<Y���>U���J-L*��{���A��ΐʠ�;�)��u��s��c��$̚3�����7
�J�<�T����R�A�J��݃�F�$b;7�]�B4G1�4^ʹ!U$�ָbMȹRT�1=��/$,2��;�.�WT����<��Xs}`Y�WԹ�E_��<�� /�[1`�G��WA�R�R	5=�D��.wO�P�+��U$2t�,"�j�y�P8#�PT�K硏�Oȕ����wp�Z��p��HS�ĳ���d�bu��-hLn�����E�����R���Q����SC��4MU��GY������xO�����5(W@*l�������G"�piKI�\��@c���T�+
�|MpSӄ)k]���� g�[rB�m�FMY�L�@�b�+��쑝;��;�%�ۣ�~ˀ|�;��b�Ӊa����Ӊ�fGE*˲�K�
�h��:��:�H�z;�ew*R���l,?��h��gf|�7�,����ϳm@A�X� < �M��T���xS�߃��~8ޥ��ưhA�oN&6���9[��c��*��~�(4�
Տ��E�� 7��ȹ��d��}+�.T�G90��"�Η�g��bެ�����@�K|}�����q�PR�~�Iz��P��qAW�����@> ~�@�<�F��qf���c�1��zJ2�����(9k_����:T��M��*+�C�؀7�i�g���{p�7���u�����m}���_#���$�������[V�om�� ]N�1�Z�"��"�j2�w@P�bJG�@���_���Ⱍ��<�JƇ�1��].\��rO�����Ln�?�ю$�c:Ye��07-���!՜'U=��R1D�gU�	콨n$�6?�]����~�dxRa����|�gD?��گ4b�q*���I��b�a�ͮDW���[O ���&�Hh���XaS�h��+�qV��ݵLBrd,�`)��?��ިq@��)-�+�Lg���=Hߴ��":�����<��D^�������|��~�jf/�;�-�*���)�z7��9�K΄�B4d��<p~Zݶ�~��W��V� ֧����F!�����B�g�Y\�����H�T��:�.ת`�V)Y���s� ���&a�?�0�����ԙSi�f��Ք��ы�(� ��|��*�!$��/�]>�Mо��H����2N���Is��0oL�/���cv��p�R���ޏ������:�T����om's���Y.:M��r�y�_�Gv��H D�ns>�c��9}N+k-�A������'���ե�6[����m���d��{q$�<�R��	�S��ɰݧj5��:���s��t ��
�e��\����j��s7�����Lyc?�<�XсP�,|���Ըp����ӽ:�+��Mxx��񕒖+����@`�̀->����� �;�u�t�W���!���	�k����x�QRp�j�S�[�zuR��N�M�h���X.��M���݅�B�
���89�0�b��%x
Wb���isI��u+�Y����K=t�i�_��@�f�#:|�fy�DS��-�p�s�'H�/�.�i�E%�s��̈́߿{W���r�'U<�_���s��G�s殾kʥ\CB�yH@`S�j7͓Zuv*�_y�W�DB*����q�)x������^�Jnsp�--F4=�	Npq�';�N���vA��.��9�I���q·���G�Bb����
 ��!]@�=tb�6�6�{�(jF3��aS^w@�i���m�Bu�g|��vd�����S�p�}��M����RB��l��Yv��u���g*���}�[)�d37D֚b-�|�g��k�y5�����Y��S�5t�Sp��� mK�����7�'8���$�DׇG�58:�,�d��A����i)�Z��6>~~U���Z��ДDn"\ƄC�3��\�`܇6�[-)��V{���x��[ȵ�|���h;AY��Q(e�N�P�cQ{ڿO>,$��R.4`졏���i0�0����1+9��kI� k��-9&C��R�ڡ������3��,%��~��
-����0t�0���4檵^��lu���2m����4j�ܬ�@����l-w}��#��K�{���B�3��U�JH()�T�K�,kA};�ph�!�=kzl>�l�$���_�h��l���Ef3���>�� �}�ǲ�WA���`��qg0��9�]Rnl9�\����&d�|�O����c�����]3�4���Q�
W2%_#,����jʌr��M��W�(}�G /{�E�*��Ђ�[|�c}�^�����k�����1 �x{"U�Χ-?�蘋c��v���a��m���=�GT��Sr4X�0�6�gS�JiK�ԓa�#�!x9b�&0R�XZ~ sZ��.�����X}Q_%<g���ͦ��N�R�C9u=׸�H���a�toME�ip�b-���@��e�d3+0��c�62">u���^TW�6Z�>7MY$��Hxh*x t���Ti����#����ϋí��M����71	�A��h���|n��eN�1�6�-A�vN,�CQ�����e�������b��B�=,�YP+�a	+h�1�.�{_M�����ؤ1��ں�<� ��dn|��A���!L:oU��;�	��y
w�H�����'��.�x�OGď Aqm���*z<B�Ѥ�1�+���H�)sHL^�^~ߥO��a��	�͊�=�V^W�7�֕(xjy� �]�U���Y�9�1 )�BO4�m�2=�8��&(8�xB�>�,���N��G�8�4���Fz3Y#�`�n�-t<@�jR�U�rȗAPＡ)/]L/��5{_�W/y�����8�ַ��Jw@E�$�r�՘���8�+3�����u����s��B��x4��� ��m��ߖɌ��\ۮ�����{�OLx����v6DK�����Z��x�7�����0�爖��/⫫�C���VUλ}=���bx��q}��" q$�=x���2_2��d8X�lq�[�fS��HO����3y?��f�ː��սz�,��:���]���Y�3r1|��;i�=ف`����-*L�}�u�k+V���7F{"��� ���'ɎT��AS-�C�|#Mz���/q<���TĊ��z;m�8��Y�����/��dB�hY�Fx�ܒ��;��w
�,�g[~���)��<�d
�Y|�U�Y�}�K4ay[�5���irh�y���R��}�����"xo#'u�!Y��ԩ�h}�x�Ѵ/{.���r�>fp�j�
>�.�f�ͨ���3�����U\�`ØJ!l%�~�'#%�pUB>l�@��Z����o���)�`b�13T凭��d��՟Asۀ�XM�$g�o��cN��44<t�'K�cIu�n�P	�J�����h8�H,���f�;����k�YY�`��Ci�V�%{�9˺$�����0μ&o��ۻ���Yb�'���O��7��@ݬ�g�>zzC����{1���d�1�J��eO��H��F�A-����f����GZ!c����x	��`*t�ܞ��\�懪_��o���I����+lI�*��7l
Ӳ�o[u8�!Ȱݾ�ٺSWQ��<�~&^k��|���8���!�R�p�r����a��U��n��$��^u
H�~[���*~eDVs�q'� �&�P����L�W����4��ѱ�x�"@.}^7�'� ���N�p0^�����5��Q��m��dԧ�*�Tb���R�x�>�$:�眮��Gu�"�]��a�+�uc��@�%�㩉^���pB���%�]��{�w
s`�����mQ�+y!���f�[k$Z���A-���v��7�.��R��4}z���ǋj,u��/�1ĩ}����2���(�BW� ��q���q���6��<�KQ�h���aX����e�9��>YF���1BG&Y��Ƴ������\�-�"���j���"���=���=�"Fq�h��?+5�����!�zA��&8p��T-�j�:gf)!�r+R�D�F$H+�&���Wx+�"��DHN�/;�&�qS;�camPL
?8�>:;}�zD��o�B*�e��b�=�e��w��=�Se*/gM8�'����z�S��.�$�oj`#�O�7�2��(}t�ӜK�9���_���ﵣç����0
](<�x�|O%"��:	`w�垵 '�x$�S�u��i��h~���\�G�׌�=�:���_=KoK���
(?�9�Փ6p�/t~h�������4TKrS����:)ɹ�R2�Y��0���[�E�ȿS-��h��\�Dt6��tL�=3�P��W�>B'W�T�Fc�l#]������h����c�l�x�M �6�@{��\��k�`�� �\���g3���&`:�����\��:ɏ[w��� 5�o�$�ATվi��)�Ѭ��V^��"p�`��������l��m�s��v���]a�k�4r)����=0�$}���ʪ<���Jܐe�I�S4zD1�����E��;�	�b�`�f�wGv� �d�H�y/� /&�q��Z7���Xr�*��:�zݱ�J��>h�e�npFN���T��gojCً.�=���{�2מq�+\z���]B�;����?��A�{j�r������Ŵ�.��ߝz�����A�t�J�	r��0~�>��J2n��*O������!h���+F(�yIN�V��a���Oi�2��v%F?#��"�p��e����C~�=�^�j<'��v��w(P8��#7<o�)�R������@�v�w��C��܍"�6~R�Ҧ��/Í�?Ws��t4]���Q\��p�B66'{��ۏN��! ���U�/�v$��|A���u<Ҁ� 1���'��#M�5VM{T��R!����iLc)1��@zd�-��(���l�<#���B�Z������F�f[�}��q�y��d�.\�C���͵�#��g)/[eR/��7��K�d�v\�V�� '*9��?[��d��VIOt/OV�TS���&�|r?p�w����[�	?�+��E�LOHh�ꖢ'��ؿ��IÈզ���XYG ̛JX�˕�nٚ�a�۔|P3��R{!����
Y\��mi�)�������fz�]�PE�����@��J�c$b��-�-�i����JN���)H;�!5� �K!q�Ů������W,��UƽPw�)cҗI���[���F���� ����5k�,�ɦ�qm��W�Ǹnf���i[/�����!�����dE���\��o��_����t��:;��x"�1,a�#��_�H�9�-
�s�ZL�9hHv}<�n��8T���9j	��)6�z��b���N��R�G�Ŵ��BE��0�{��.M	||�>��-D��uö���J}@�l�5r�ޥ�A}^?��Cc�E�b�"��a	ا��虢�m��*ģ�#� 	R�9P�ʸ�j�B%��sFJΖ��Z���;Q�j��;��w�t�{������k��A��|xG`��.$�d�%��rup8' [0�f�fR��l}	�&�*�V���f�
m�%Xk�ceu[�;�EtV��"�Iw'k�&E�;�r������)��ة��5��X��?�
��#1�-��R�G���$�ʄ躸S�P�N��V
ʣ�)w���>����3�B��Mj����N{[�5�\����0���#�S�,�ս���u�R~��r�>�x��/��zB��S%�{�P{AŪg����V"�ݡ�����&���6���~��e�
�#��U-F���
LfԸ�@������rZ�+���z�~I��#z��:נ�����T���be�C;#־���pSe2�M�Մ��s7ւ�$/� ���=ŔV<M�ׯ��Pd68UO~�g4zӭru�m�?��;�N����T�ѭ�Q�c�G����K>��j�>U��G�C�&}qᐜ�Q~������&���{�k�mF�}4�ُ�P`��	����7Xt[�Y�/�.��u-!K�@s����0E+Z�-9P�A���|V;`�f�[�v���L �2��wްS�|,�<�L1�Ú
Z����bq�<;���>�/�n6U�u�i�s���+���Bg�^0��k���t �sG,	~�� /��f�	���(6�����;ڎv��C)�%�O�,�.����B���hIg\�-e[QS��X<6�Oh��h-o���v<Z!sd�ۈ��m%B��zR݋��K��k>� V�9l\�����f��_�
����E�C��_�K���g�I�@;�[����j�,:��2�T��TJ�����׬|��&g�����W�ﵖr!ͯ�ٶ�I1��gʽ�mȈʢ�W����@Tϔ��XF|�6����p���a��v7�@%�(WaTg�L���z�=.e�2�����G�*��!�$1�[������*m��̉J`�e&����h��c8�N�?F�&ɭ��R��R!�����A�G�;�fH�����^��N�[1"���
��i�<����+��q\�C�	O����=s��+<�q�TRR�U�m��������ѱ0�1ƓP�h�	5@%ʄ�mq����=�W@>�L���)<��p�+��z����PsL�Yf����C����'ҴT�aE�>K�p�;��SR�-���"����"`Q�0���to]�]�x�!տ%�������*^i���YB�G��Y�
ش�MB ��yyy�	���5[���SR)^V+�)�+�V��u�}��Wq|�j����QI�d�ƽ[Ɠ�GI���vc��uJ��&�K�PI�����>��Dc47lo�2�M��8,�y�B���3��{���5Pi��_�mƣ�A+1O0���$������5����i��TL�mr�O�nml�Y���yݽ��*ȡ4�v���r'�S~����5������խ�>���N8�jG��EB�M̳Ia�+|�8'��cG�a�./�Z��%�ԉL�<�FHS`^���~�.��%�l~��R���ZfJ1���8�_0�)Ĵ���TxNJs�[� e/T�|x_VO��x��B�g��f���%\k�(ʘ#;�o��~< �*A��Ag�����U'�6>2�Ҏ�[�_K�y���U���fcy��$7W8杢�#:˄;�Ⱥ�5�k���Q�x��8���̕�K�(����6i�<���9Wy#e�����*���
�2��"�u}�i�J����8^8d<���E)�2�k��`�-�&De�+�F��[h�Я�V��B�0(���l�\�c�4PBW�$g��!4��A:n���h��oG�TH��O	þ��(ami�B��j��_tyo�\aÔk���>����z��4e�̨`�bO�P�V29��A-C�P�Z5��ӊ�N�/4��]��~���7�Mp������y��˲�uT74���ѫ\���Ut�v�c�&#9a�ҍ�J�	�%��Ɍue����J�B��!�͙~%.֪ɔ�X�C��GRU;r?]$6U}�����=���j��F��X�,�/�F�L�A����1(uh�7	ÂX.�h+�]7��EVx�:!*�2���%,�q��A~+zQ�fL���j�8�0k����]bR��k��NC��J��?fb/�Z���$d4{���TΡ�&��v�)I��,��ޑ2���
�#{W�3�Q�����w*$m�p!V{k���9��3��Y�`�BO��˫�����9�4��(<���0�\�1���������EYS�n-1U/ԩZ 7���Z�b*5��Z-((O�	������	�J�Ȇ^P">�����E��#P�8�r9'����x�"��N�K��L��Nh�N�SG��ۦ�^�W�;㍳��C��EHƍ���� ���zV�K��*{���9xmҏ�7J���Y�hΪ�FNe�F�u�7�GcKU��pm�ś���4Pݎg2������I_�`W@�Ȉ�LPs(c�-D��u,� m������Y�s�i%j������~H8��wO�H���jo�Q�k�p嬶����ҫ��D�۴�+�d۠�T#!{\�;�,А��R����A��0+��4ٗ.�B^�k�&U�a�؋������:bgl�j���|=�R%�PH7v�h�]��P�NG[���{r�^$=�A�E�6I�Uo�8MR��$4}���QD�0K|�N���f��[��5�rYZ0KU?TjY�x�������V�v��E��pf�����}/�՞�!����?�HF�nR��|��׆�Iu�o�}'H�90�ߑi�m忉	\�������}.�ȼ*��^�����uOo��Y/��l�R�չ9����_��t_�M�2������5��u���?�y>�.�%���U�����ey{��� � {M�����m�u׻���y���~Ik�!����;F�����d)��@Ԅ��.��_7c��\�5�{������E��bP��u��*l�V7�`�~�K�_�Z�2�)���k��_)�
&|����p�#�2��u� H,��顚��<�٠�jaVY [_��z��G�)wY��>gj�ﭚóM� س�c� oZzh����c���n�A]U��ڈ\��1B�D���=?��l��}GaOa%ZU1��Q��Q�ߑ�k�N�Z�M)�q��P# �~�N[�n/U�.7�+���g�Z���� $2$SA<�z����1��{a'!k�Pn�#��Q�֖����0�ۊ��S��]G�ts�����""\�O.J�)俇oᵙ^ru�R�]�d��|L���OȈC�-�`�L'*���ƅZ�6�� �W�R�S}�i��ahU/���WK���@��D��ٶ�񕰎�I|eC�+R��3u��h��
?o�o��i�K՟����Z[m��re�Y�|����i9f���� eRē�y�� ����U-��5��cA�}sjɓ�t H�Μ��f&�Ӽ٤K߱���"�U���Y<=f�Y�Ǉ�� �%2�>����rb��C��Wh�Zh������>���+�Q7��k]�'R��Bu�ؼ�CgU�\�T7*��ҤE��� ��X���a�16�=���)-�j�8��6i]�F��8�����B�3h��f����s�ߦ�ԡ��mM���-{h&Xd�yX�P�i�+�O�4�юYh�<�U��sQ�<K[�r��iv���-�s��uOO��Di��(����>�I�ɳ�V�!;&�%��0���Iy0�gW?!V���B��﹪X�oL5�s��f�R;��M���LK��ٸ1���4-FQNp��$��/8زr��S��s"��6�Z��)u��5�6,V�ڂ�@��G�R�W)���!s41{���bc�^֘�OJa����#y~�=v-��S�ˉ$���e�U�!G!J��C��R�V�E��d��|a�3ً&փ���o��3.jѷ��&�'��f�(���^%�P,��O��K�q's.�'oI�M�:7��^���p�ʳ,r�c�[���t۴��3�xQ��T5�&{1 ���q�Ǧ��=�GѪG����q#3�i��� ��������۠U7wF��np�%fZ�����з��rv�P��w�޸Llo�^����������������1�);CGQ���M����rz�[@�M���O�����*�~,�k9����w����A1G�`p��r�-�$�`&�C�{�[���Y~�y��e����RZ1A����u^M��	X��>�h��峝��t��=���iL�^��sY���1"6��R��9��(�ϒ���Q�5�E�_͋~�T��0�醦%bU4�횙��ʃ�s} (+�A����o�Ğ��,(q[v�.Q{3�^�O���ׯ��n�����r�{�\��Y%�1Mʾ~e��
�<
C��u�/J��iT[���_8G���-I0Y�a���Nhv��^��"�t���ҧ!w�)�NVD6�7Y�L��cɖ��f�&U֬�]�eKwTY?
GYR�+#�I��y�|J���BA�;ef*m�"�(�6�T=�
p �24�b�>΄�0`�L�[�|��R�OR�Ո�#� H��H���u{[S��	�QܤҲ|	J,mj�4J��<o6��K60o�i�~�+{�Ɠ��54T=�u��o��sõ��b�ܖ�&q��|���'�7�v�T6Ɠ�\���T����Fa-q���0�D⾫�[��hk$�9����Ё�}ɧ&�e�����A �$�k�C%�tČ�9]΂�bΐH�X�|����#T�Xh��1O5qJ�uɌ�Z
-���^�����7�r�ǇP7���'��%���vzbƲ|Y�����2�����ԁ2+�������*��}a��{+�4_ �d}נ�o��MP�=�!�'�|��߹�]����&
�C�b�#�B��G��|j�[cc�G�C��uF"�fq͝534l�����)un	��p�����P4�kwd���0i�P��3z�r��M�z��;L�s�u�[4s�.�c62/�X#����*�x�;�I��a�\�����5���qզ1�S��2|b����&�V{P���N-ԅY_�y�J޳ e������$J-�o�hF=�D����}�p|t��Q�h���}WxL�?��f��3�G�U���[ƇZ� ��)��?��4P�Ӛ�Չ��(H�$1ᙳ�.�\#�Vݸ�9�:�2+���'�?m����,x��t�x��+��\�ɉP)��^z�϶��ْ�0�q�iI��֎-�Whe��zK���i{��ֱ��],�����/�#�������ʤ�4��By[���;�uq��>ж|q�~���rd2��%_���5/R����1�������N@E;�D,�]'�ݣRL�Qc���LG!rIyh�����LJ�v���
v{2�H�w��CĀ��X�UȌN�����wxi��;��(����������w�0��	�u�-�{�s����c����'d�޵۝G��n@�x�����������&"��d�����=v�2,waQfD�^�f�]���ߔS��tF�<bM3�-�,Hہثi����~1�z)���a]�9|��������퉕0J�,>WR-�=��ΛҲ�������Ϲs�-6^�`����pӏ�}-bX6`m?�i���@Gwܝz�~F��{�>0��Ll��{G��|xS�vUl��1�h���U�b�RI�R��۩�u~y��?��1W���jW@/c�b�Ga�т���9l�ܩyMܽ�eֶ ϣv�ku�ڑ_���햆������D�3�l�x�â��˅Ģ�C�F6�:������	�)&ʡ������U���t���hEx���ᑉ_[�IF8Ӫ_R%V7�����,�ЃƤ �-U��LZ�P�� O�g}<�5��1��X���ܺ�߻0�_6��ɶh&1&`x��2Dp�����8�(����aFĮ�
��?����Af(��֣�{���\����:C����s$ʄ�FU��P�O����B�#�b����k"�ciz����q"�R�g�]&�t��{<U����+�@��
<�	��f2� ���M"����= �'8�:׃��iů�B"�W)���r�}Q3�p�z����P�~FK�ò��-� �m�{��L�g�<�'��]�~�m�ͦK�L��<�&��Y���8��d-'�V���9�aG
䬑�ĥ܍m��EЖ�-��uʌ��	D>��J�p.��m����Nrzԧ?��J�,9���A�_Lpb Ҋ�6�
�{'���H�~�����0�θ�� ��d}���}&�UîG���'�zgW^���<]2�eޗ,�8Phۘ�J~I5�[R����Ұ'���I�"����2CГ.)F����Բ�m#��I�Ыbɘ��~���C>,y-�}I�v����s��Yw@��]��	�k�5������U ~p6�Q��$��9j�㾢��/����g��)i�a�P	�Ҁ� BP3 ����r��8�WSΜ�*�����n�P4C�i�-��
�cLE�AP�7�3�t;K����N����3�i���[s@[����Ac�)����+�{V�$^WTR�6FN@^1�BU�.�	��V?������2�T��۞z�ѥ߯�C��k�a�nW!ib�<�x2��zuk{w�'���\�����<=�JV��"��!$��
���L_#T�[y�^�� 'x���۪�귞/�	cx�q��́r�"S����Ik(�q�J�Ma,��Y~,�|��d��m0jٙt1�i4O�^�������Z�'lI�So5G�	<���'[0~o�G_):.+	���γ8n�&�gM��2S�W����7o��B�ǃ_o1+Wl<
V��'|�����t��;x7uE���L��ʞ��(a:��4i��i�_����c(7��=!�B���.ZS�t�2)�>a��|�)&��+(UWx�k���Y�]MuwaTii��P��7�{Q��Ǔ[ ��eW��$ʾ�x.�Y�^�\����D�C���yu��z�\	?fD�#jA��Ք#�S~���Ԍ���Iӫ)�9��?�WQŤ�
��~�j*�
%EL
G�7�4�q~ ���ؕ��Í���9��a�G埶�h8�zo��a��AI٦��50߈I"�+��?�E�#=�?T�0�\V�z��+���M�Ӧi�ɇ	�hd��S	lh9K����_gc2g1\x��_�|��.�C�O^^�Ǣ���rM�ڎn��c�$�9]��Kޢ���$�LE���{�H[�