-- DOC_Monitor.vhd

-- Generated using ACDS version 14.0 200 at 2015.05.08.14:44:54

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DOC_Monitor is
	port (
		in_port_to_the_IO_IN_Buttons   : in  std_logic_vector(3 downto 0)  := (others => '0'); -- io_in_buttons_external_connection.export
		pio_pfc_in_port                : in  std_logic_vector(1 downto 0)  := (others => '0'); --                           pio_pfc.in_port
		pio_pfc_out_port               : out std_logic_vector(1 downto 0);                     --                                  .out_port
		dc_link_sync_dat               : in  std_logic                     := '0';             --                           dc_link.sync_dat
		dc_link_dc_link_enable         : in  std_logic                     := '0';             --                                  .dc_link_enable
		dc_link_overvoltage            : out std_logic;                                        --                                  .overvoltage
		dc_link_undervoltage           : out std_logic;                                        --                                  .undervoltage
		dc_link_chopper                : out std_logic;                                        --                                  .chopper
		dc_link_p_sync_dat             : in  std_logic                     := '0';             --                         dc_link_p.sync_dat
		dc_link_p_dc_link_enable       : in  std_logic                     := '0';             --                                  .dc_link_enable
		dc_link_p_overvoltage          : out std_logic;                                        --                                  .overvoltage
		dc_link_p_undervoltage         : out std_logic;                                        --                                  .undervoltage
		dc_link_p_chopper              : out std_logic;                                        --                                  .chopper
		clk_adc_in_clk                 : in  std_logic                     := '0';             --                        clk_adc_in.clk
		avs_periph_slave_waitrequest   : out std_logic;                                        --                  avs_periph_slave.waitrequest
		avs_periph_slave_readdata      : out std_logic_vector(31 downto 0);                    --                                  .readdata
		avs_periph_slave_readdatavalid : out std_logic;                                        --                                  .readdatavalid
		avs_periph_slave_burstcount    : in  std_logic_vector(0 downto 0)  := (others => '0'); --                                  .burstcount
		avs_periph_slave_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --                                  .writedata
		avs_periph_slave_address       : in  std_logic_vector(11 downto 0) := (others => '0'); --                                  .address
		avs_periph_slave_write         : in  std_logic                     := '0';             --                                  .write
		avs_periph_slave_read          : in  std_logic                     := '0';             --                                  .read
		avs_periph_slave_byteenable    : in  std_logic_vector(3 downto 0)  := (others => '0'); --                                  .byteenable
		avs_periph_slave_debugaccess   : in  std_logic                     := '0';             --                                  .debugaccess
		clk_80_clk                     : in  std_logic                     := '0';             --                            clk_80.clk
		reset_80_reset_n               : in  std_logic                     := '0';             --                          reset_80.reset_n
		clk_50_clk                     : in  std_logic                     := '0';             --                            clk_50.clk
		reset_50_reset_n               : in  std_logic                     := '0'              --                          reset_50.reset_n
	);
end entity DOC_Monitor;

architecture rtl of DOC_Monitor is
	component DOC_Monitor_IO_IN_Buttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component DOC_Monitor_IO_IN_Buttons;

	component altera_avalon_mm_clock_crossing_bridge is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			HDL_ADDR_WIDTH      : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(11 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component altera_avalon_mm_clock_crossing_bridge;

	component ssg_emb_dc_ballast is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			avs_write_n    : in  std_logic                     := 'X';             -- write_n
			avs_read_n     : in  std_logic                     := 'X';             -- read_n
			avs_address    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avs_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			reset_n        : in  std_logic                     := 'X';             -- reset_n
			sync_dat       : in  std_logic                     := 'X';             -- export
			dc_link_enable : in  std_logic                     := 'X';             -- export
			overvoltage    : out std_logic;                                        -- export
			undervoltage   : out std_logic;                                        -- export
			chopper        : out std_logic;                                        -- export
			clk_adc        : in  std_logic                     := 'X'              -- clk
		);
	end component ssg_emb_dc_ballast;

	component DOC_Monitor_pio_pfc is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component DOC_Monitor_pio_pfc;

	component DOC_Monitor_sysid_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component DOC_Monitor_sysid_0;

	component DOC_Monitor_mm_interconnect_0 is
		port (
			clk_int_50_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			clock_crossing_m0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			clock_crossing_m0_address                           : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			clock_crossing_m0_waitrequest                       : out std_logic;                                        -- waitrequest
			clock_crossing_m0_burstcount                        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			clock_crossing_m0_byteenable                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clock_crossing_m0_read                              : in  std_logic                     := 'X';             -- read
			clock_crossing_m0_readdata                          : out std_logic_vector(31 downto 0);                    -- readdata
			clock_crossing_m0_readdatavalid                     : out std_logic;                                        -- readdatavalid
			clock_crossing_m0_write                             : in  std_logic                     := 'X';             -- write
			clock_crossing_m0_writedata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clock_crossing_m0_debugaccess                       : in  std_logic                     := 'X';             -- debugaccess
			DOC_DC_Link_avalon_slave_0_address                  : out std_logic_vector(3 downto 0);                     -- address
			DOC_DC_Link_avalon_slave_0_write                    : out std_logic;                                        -- write
			DOC_DC_Link_avalon_slave_0_read                     : out std_logic;                                        -- read
			DOC_DC_Link_avalon_slave_0_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DOC_DC_Link_avalon_slave_0_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			DOC_DC_Link_P_avalon_slave_0_address                : out std_logic_vector(3 downto 0);                     -- address
			DOC_DC_Link_P_avalon_slave_0_write                  : out std_logic;                                        -- write
			DOC_DC_Link_P_avalon_slave_0_read                   : out std_logic;                                        -- read
			DOC_DC_Link_P_avalon_slave_0_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DOC_DC_Link_P_avalon_slave_0_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			IO_IN_Buttons_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			IO_IN_Buttons_s1_write                              : out std_logic;                                        -- write
			IO_IN_Buttons_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			IO_IN_Buttons_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			IO_IN_Buttons_s1_chipselect                         : out std_logic;                                        -- chipselect
			pio_pfc_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			pio_pfc_s1_write                                    : out std_logic;                                        -- write
			pio_pfc_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_pfc_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			pio_pfc_s1_chipselect                               : out std_logic;                                        -- chipselect
			sysid_0_control_slave_address                       : out std_logic_vector(0 downto 0);                     -- address
			sysid_0_control_slave_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component DOC_Monitor_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal clock_crossing_m0_burstcount                                   : std_logic_vector(0 downto 0);  -- clock_crossing:m0_burstcount -> mm_interconnect_0:clock_crossing_m0_burstcount
	signal clock_crossing_m0_waitrequest                                  : std_logic;                     -- mm_interconnect_0:clock_crossing_m0_waitrequest -> clock_crossing:m0_waitrequest
	signal clock_crossing_m0_address                                      : std_logic_vector(11 downto 0); -- clock_crossing:m0_address -> mm_interconnect_0:clock_crossing_m0_address
	signal clock_crossing_m0_writedata                                    : std_logic_vector(31 downto 0); -- clock_crossing:m0_writedata -> mm_interconnect_0:clock_crossing_m0_writedata
	signal clock_crossing_m0_write                                        : std_logic;                     -- clock_crossing:m0_write -> mm_interconnect_0:clock_crossing_m0_write
	signal clock_crossing_m0_read                                         : std_logic;                     -- clock_crossing:m0_read -> mm_interconnect_0:clock_crossing_m0_read
	signal clock_crossing_m0_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:clock_crossing_m0_readdata -> clock_crossing:m0_readdata
	signal clock_crossing_m0_debugaccess                                  : std_logic;                     -- clock_crossing:m0_debugaccess -> mm_interconnect_0:clock_crossing_m0_debugaccess
	signal clock_crossing_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- clock_crossing:m0_byteenable -> mm_interconnect_0:clock_crossing_m0_byteenable
	signal clock_crossing_m0_readdatavalid                                : std_logic;                     -- mm_interconnect_0:clock_crossing_m0_readdatavalid -> clock_crossing:m0_readdatavalid
	signal mm_interconnect_0_io_in_buttons_s1_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:IO_IN_Buttons_s1_writedata -> IO_IN_Buttons:writedata
	signal mm_interconnect_0_io_in_buttons_s1_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:IO_IN_Buttons_s1_address -> IO_IN_Buttons:address
	signal mm_interconnect_0_io_in_buttons_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:IO_IN_Buttons_s1_chipselect -> IO_IN_Buttons:chipselect
	signal mm_interconnect_0_io_in_buttons_s1_write                       : std_logic;                     -- mm_interconnect_0:IO_IN_Buttons_s1_write -> mm_interconnect_0_io_in_buttons_s1_write:in
	signal mm_interconnect_0_io_in_buttons_s1_readdata                    : std_logic_vector(31 downto 0); -- IO_IN_Buttons:readdata -> mm_interconnect_0:IO_IN_Buttons_s1_readdata
	signal mm_interconnect_0_doc_dc_link_avalon_slave_0_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:DOC_DC_Link_avalon_slave_0_writedata -> DOC_DC_Link:avs_writedata
	signal mm_interconnect_0_doc_dc_link_avalon_slave_0_address           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:DOC_DC_Link_avalon_slave_0_address -> DOC_DC_Link:avs_address
	signal mm_interconnect_0_doc_dc_link_avalon_slave_0_write             : std_logic;                     -- mm_interconnect_0:DOC_DC_Link_avalon_slave_0_write -> mm_interconnect_0_doc_dc_link_avalon_slave_0_write:in
	signal mm_interconnect_0_doc_dc_link_avalon_slave_0_read              : std_logic;                     -- mm_interconnect_0:DOC_DC_Link_avalon_slave_0_read -> mm_interconnect_0_doc_dc_link_avalon_slave_0_read:in
	signal mm_interconnect_0_doc_dc_link_avalon_slave_0_readdata          : std_logic_vector(31 downto 0); -- DOC_DC_Link:avs_readdata -> mm_interconnect_0:DOC_DC_Link_avalon_slave_0_readdata
	signal mm_interconnect_0_doc_dc_link_p_avalon_slave_0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:DOC_DC_Link_P_avalon_slave_0_writedata -> DOC_DC_Link_P:avs_writedata
	signal mm_interconnect_0_doc_dc_link_p_avalon_slave_0_address         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:DOC_DC_Link_P_avalon_slave_0_address -> DOC_DC_Link_P:avs_address
	signal mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write           : std_logic;                     -- mm_interconnect_0:DOC_DC_Link_P_avalon_slave_0_write -> mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write:in
	signal mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read            : std_logic;                     -- mm_interconnect_0:DOC_DC_Link_P_avalon_slave_0_read -> mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read:in
	signal mm_interconnect_0_doc_dc_link_p_avalon_slave_0_readdata        : std_logic_vector(31 downto 0); -- DOC_DC_Link_P:avs_readdata -> mm_interconnect_0:DOC_DC_Link_P_avalon_slave_0_readdata
	signal mm_interconnect_0_pio_pfc_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_pfc_s1_writedata -> pio_pfc:writedata
	signal mm_interconnect_0_pio_pfc_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_pfc_s1_address -> pio_pfc:address
	signal mm_interconnect_0_pio_pfc_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:pio_pfc_s1_chipselect -> pio_pfc:chipselect
	signal mm_interconnect_0_pio_pfc_s1_write                             : std_logic;                     -- mm_interconnect_0:pio_pfc_s1_write -> mm_interconnect_0_pio_pfc_s1_write:in
	signal mm_interconnect_0_pio_pfc_s1_readdata                          : std_logic_vector(31 downto 0); -- pio_pfc:readdata -> mm_interconnect_0:pio_pfc_s1_readdata
	signal mm_interconnect_0_sysid_0_control_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_0_control_slave_address -> sysid_0:address
	signal mm_interconnect_0_sysid_0_control_slave_readdata               : std_logic_vector(31 downto 0); -- sysid_0:readdata -> mm_interconnect_0:sysid_0_control_slave_readdata
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [clock_crossing:m0_reset, mm_interconnect_0:clock_crossing_m0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                             : std_logic;                     -- rst_controller_001:reset_out -> clock_crossing:s0_reset
	signal reset_80_reset_n_ports_inv                                     : std_logic;                     -- reset_80_reset_n:inv -> rst_controller_001:reset_in0
	signal reset_50_reset_n_ports_inv                                     : std_logic;                     -- reset_50_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_io_in_buttons_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_0_io_in_buttons_s1_write:inv -> IO_IN_Buttons:write_n
	signal mm_interconnect_0_doc_dc_link_avalon_slave_0_write_ports_inv   : std_logic;                     -- mm_interconnect_0_doc_dc_link_avalon_slave_0_write:inv -> DOC_DC_Link:avs_write_n
	signal mm_interconnect_0_doc_dc_link_avalon_slave_0_read_ports_inv    : std_logic;                     -- mm_interconnect_0_doc_dc_link_avalon_slave_0_read:inv -> DOC_DC_Link:avs_read_n
	signal mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write_ports_inv : std_logic;                     -- mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write:inv -> DOC_DC_Link_P:avs_write_n
	signal mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read_ports_inv  : std_logic;                     -- mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read:inv -> DOC_DC_Link_P:avs_read_n
	signal mm_interconnect_0_pio_pfc_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_pio_pfc_s1_write:inv -> pio_pfc:write_n
	signal rst_controller_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_reset_out_reset:inv -> [DOC_DC_Link:reset_n, DOC_DC_Link_P:reset_n, IO_IN_Buttons:reset_n, pio_pfc:reset_n, sysid_0:reset_n]

begin

	io_in_buttons : component DOC_Monitor_IO_IN_Buttons
		port map (
			clk        => clk_50_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_io_in_buttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_io_in_buttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_io_in_buttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_io_in_buttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_io_in_buttons_s1_readdata,        --                    .readdata
			in_port    => in_port_to_the_IO_IN_Buttons                        -- external_connection.export
		);

	clock_crossing : component altera_avalon_mm_clock_crossing_bridge
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			HDL_ADDR_WIDTH      => 12,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 2,
			RESPONSE_FIFO_DEPTH => 2,
			MASTER_SYNC_DEPTH   => 3,
			SLAVE_SYNC_DEPTH    => 3
		)
		port map (
			m0_clk           => clk_50_clk,                         --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,     -- m0_reset.reset
			s0_clk           => clk_80_clk,                         --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset, -- s0_reset.reset
			s0_waitrequest   => avs_periph_slave_waitrequest,       --       s0.waitrequest
			s0_readdata      => avs_periph_slave_readdata,          --         .readdata
			s0_readdatavalid => avs_periph_slave_readdatavalid,     --         .readdatavalid
			s0_burstcount    => avs_periph_slave_burstcount,        --         .burstcount
			s0_writedata     => avs_periph_slave_writedata,         --         .writedata
			s0_address       => avs_periph_slave_address,           --         .address
			s0_write         => avs_periph_slave_write,             --         .write
			s0_read          => avs_periph_slave_read,              --         .read
			s0_byteenable    => avs_periph_slave_byteenable,        --         .byteenable
			s0_debugaccess   => avs_periph_slave_debugaccess,       --         .debugaccess
			m0_waitrequest   => clock_crossing_m0_waitrequest,      --       m0.waitrequest
			m0_readdata      => clock_crossing_m0_readdata,         --         .readdata
			m0_readdatavalid => clock_crossing_m0_readdatavalid,    --         .readdatavalid
			m0_burstcount    => clock_crossing_m0_burstcount,       --         .burstcount
			m0_writedata     => clock_crossing_m0_writedata,        --         .writedata
			m0_address       => clock_crossing_m0_address,          --         .address
			m0_write         => clock_crossing_m0_write,            --         .write
			m0_read          => clock_crossing_m0_read,             --         .read
			m0_byteenable    => clock_crossing_m0_byteenable,       --         .byteenable
			m0_debugaccess   => clock_crossing_m0_debugaccess       --         .debugaccess
		);

	doc_dc_link : component ssg_emb_dc_ballast
		port map (
			clk            => clk_50_clk,                                                   --          clock.clk
			avs_write_n    => mm_interconnect_0_doc_dc_link_avalon_slave_0_write_ports_inv, -- avalon_slave_0.write_n
			avs_read_n     => mm_interconnect_0_doc_dc_link_avalon_slave_0_read_ports_inv,  --               .read_n
			avs_address    => mm_interconnect_0_doc_dc_link_avalon_slave_0_address,         --               .address
			avs_writedata  => mm_interconnect_0_doc_dc_link_avalon_slave_0_writedata,       --               .writedata
			avs_readdata   => mm_interconnect_0_doc_dc_link_avalon_slave_0_readdata,        --               .readdata
			reset_n        => rst_controller_reset_out_reset_ports_inv,                     --          reset.reset_n
			sync_dat       => dc_link_sync_dat,                                             --         status.export
			dc_link_enable => dc_link_dc_link_enable,                                       --               .export
			overvoltage    => dc_link_overvoltage,                                          --               .export
			undervoltage   => dc_link_undervoltage,                                         --               .export
			chopper        => dc_link_chopper,                                              --               .export
			clk_adc        => clk_adc_in_clk                                                --      clock_adc.clk
		);

	doc_dc_link_p : component ssg_emb_dc_ballast
		port map (
			clk            => clk_50_clk,                                                     --          clock.clk
			avs_write_n    => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write_ports_inv, -- avalon_slave_0.write_n
			avs_read_n     => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read_ports_inv,  --               .read_n
			avs_address    => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_address,         --               .address
			avs_writedata  => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_writedata,       --               .writedata
			avs_readdata   => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_readdata,        --               .readdata
			reset_n        => rst_controller_reset_out_reset_ports_inv,                       --          reset.reset_n
			sync_dat       => dc_link_p_sync_dat,                                             --         status.export
			dc_link_enable => dc_link_p_dc_link_enable,                                       --               .export
			overvoltage    => dc_link_p_overvoltage,                                          --               .export
			undervoltage   => dc_link_p_undervoltage,                                         --               .export
			chopper        => dc_link_p_chopper,                                              --               .export
			clk_adc        => clk_adc_in_clk                                                  --      clock_adc.clk
		);

	pio_pfc : component DOC_Monitor_pio_pfc
		port map (
			clk        => clk_50_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pio_pfc_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_pfc_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_pfc_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_pfc_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_pfc_s1_readdata,        --                    .readdata
			in_port    => pio_pfc_in_port,                              -- external_connection.export
			out_port   => pio_pfc_out_port                              --                    .export
		);

	sysid_0 : component DOC_Monitor_sysid_0
		port map (
			clock    => clk_50_clk,                                         --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,           --         reset.reset_n
			readdata => mm_interconnect_0_sysid_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component DOC_Monitor_mm_interconnect_0
		port map (
			clk_int_50_clk_clk                                  => clk_50_clk,                                               --                                clk_int_50_clk.clk
			clock_crossing_m0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                           -- clock_crossing_m0_reset_reset_bridge_in_reset.reset
			clock_crossing_m0_address                           => clock_crossing_m0_address,                                --                             clock_crossing_m0.address
			clock_crossing_m0_waitrequest                       => clock_crossing_m0_waitrequest,                            --                                              .waitrequest
			clock_crossing_m0_burstcount                        => clock_crossing_m0_burstcount,                             --                                              .burstcount
			clock_crossing_m0_byteenable                        => clock_crossing_m0_byteenable,                             --                                              .byteenable
			clock_crossing_m0_read                              => clock_crossing_m0_read,                                   --                                              .read
			clock_crossing_m0_readdata                          => clock_crossing_m0_readdata,                               --                                              .readdata
			clock_crossing_m0_readdatavalid                     => clock_crossing_m0_readdatavalid,                          --                                              .readdatavalid
			clock_crossing_m0_write                             => clock_crossing_m0_write,                                  --                                              .write
			clock_crossing_m0_writedata                         => clock_crossing_m0_writedata,                              --                                              .writedata
			clock_crossing_m0_debugaccess                       => clock_crossing_m0_debugaccess,                            --                                              .debugaccess
			DOC_DC_Link_avalon_slave_0_address                  => mm_interconnect_0_doc_dc_link_avalon_slave_0_address,     --                    DOC_DC_Link_avalon_slave_0.address
			DOC_DC_Link_avalon_slave_0_write                    => mm_interconnect_0_doc_dc_link_avalon_slave_0_write,       --                                              .write
			DOC_DC_Link_avalon_slave_0_read                     => mm_interconnect_0_doc_dc_link_avalon_slave_0_read,        --                                              .read
			DOC_DC_Link_avalon_slave_0_readdata                 => mm_interconnect_0_doc_dc_link_avalon_slave_0_readdata,    --                                              .readdata
			DOC_DC_Link_avalon_slave_0_writedata                => mm_interconnect_0_doc_dc_link_avalon_slave_0_writedata,   --                                              .writedata
			DOC_DC_Link_P_avalon_slave_0_address                => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_address,   --                  DOC_DC_Link_P_avalon_slave_0.address
			DOC_DC_Link_P_avalon_slave_0_write                  => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write,     --                                              .write
			DOC_DC_Link_P_avalon_slave_0_read                   => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read,      --                                              .read
			DOC_DC_Link_P_avalon_slave_0_readdata               => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_readdata,  --                                              .readdata
			DOC_DC_Link_P_avalon_slave_0_writedata              => mm_interconnect_0_doc_dc_link_p_avalon_slave_0_writedata, --                                              .writedata
			IO_IN_Buttons_s1_address                            => mm_interconnect_0_io_in_buttons_s1_address,               --                              IO_IN_Buttons_s1.address
			IO_IN_Buttons_s1_write                              => mm_interconnect_0_io_in_buttons_s1_write,                 --                                              .write
			IO_IN_Buttons_s1_readdata                           => mm_interconnect_0_io_in_buttons_s1_readdata,              --                                              .readdata
			IO_IN_Buttons_s1_writedata                          => mm_interconnect_0_io_in_buttons_s1_writedata,             --                                              .writedata
			IO_IN_Buttons_s1_chipselect                         => mm_interconnect_0_io_in_buttons_s1_chipselect,            --                                              .chipselect
			pio_pfc_s1_address                                  => mm_interconnect_0_pio_pfc_s1_address,                     --                                    pio_pfc_s1.address
			pio_pfc_s1_write                                    => mm_interconnect_0_pio_pfc_s1_write,                       --                                              .write
			pio_pfc_s1_readdata                                 => mm_interconnect_0_pio_pfc_s1_readdata,                    --                                              .readdata
			pio_pfc_s1_writedata                                => mm_interconnect_0_pio_pfc_s1_writedata,                   --                                              .writedata
			pio_pfc_s1_chipselect                               => mm_interconnect_0_pio_pfc_s1_chipselect,                  --                                              .chipselect
			sysid_0_control_slave_address                       => mm_interconnect_0_sysid_0_control_slave_address,          --                         sysid_0_control_slave.address
			sysid_0_control_slave_readdata                      => mm_interconnect_0_sysid_0_control_slave_readdata          --                                              .readdata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_50_reset_n_ports_inv,     -- reset_in0.reset
			clk            => clk_50_clk,                     --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_80_reset_n_ports_inv,         -- reset_in0.reset
			clk            => clk_80_clk,                         --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_80_reset_n_ports_inv <= not reset_80_reset_n;

	reset_50_reset_n_ports_inv <= not reset_50_reset_n;

	mm_interconnect_0_io_in_buttons_s1_write_ports_inv <= not mm_interconnect_0_io_in_buttons_s1_write;

	mm_interconnect_0_doc_dc_link_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_doc_dc_link_avalon_slave_0_write;

	mm_interconnect_0_doc_dc_link_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_doc_dc_link_avalon_slave_0_read;

	mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_doc_dc_link_p_avalon_slave_0_write;

	mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_doc_dc_link_p_avalon_slave_0_read;

	mm_interconnect_0_pio_pfc_s1_write_ports_inv <= not mm_interconnect_0_pio_pfc_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of DOC_Monitor
